//
// Copyright (c) 2016 University of Cambridge All rights reserved.
//
// Author: Marco Forconesi
//
// This software was developed with the support of
// Prof. Gustavo Sutter and Prof. Sergio Lopez-Buedo and
// University of Cambridge Computer Laboratory NetFPGA team.
//
// @NETFPGA_LICENSE_HEADER_START@
//
// Licensed to NetFPGA C.I.C. (NetFPGA) under one or more
// contributor license agreements.  See the NOTICE file distributed with this
// work for additional information regarding copyright ownership.  NetFPGA
// licenses this file to you under the NetFPGA Hardware-Software License,
// Version 1.0 (the "License"); you may not use this file except in compliance
// with the License.  You may obtain a copy of the License at:
//
//   http://www.netfpga-cic.org
//
// Unless required by applicable law or agreed to in writing, Work distributed
// under the License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied.  See the License for the
// specific language governing permissions and limitations under the License.
//
// @NETFPGA_LICENSE_HEADER_END@

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

    // XGMII characters
    localparam S   = 8'hFB;
    localparam T   = 8'hFD;
    localparam E   = 8'hFE;
    localparam I   = 8'h07;

    localparam PREAMBLE_LANE0_D = {56'hD5555555555555, S};
    localparam PREAMBLE_LANE0_C = 8'h01;

    localparam PREAMBLE_LANE4_D = {24'h555555, S, {4{I}}};
    localparam PREAMBLE_LANE4_C = 8'h1F;

    localparam PREAMBLE_LANE4_END_D = 32'hD5555555;
    localparam PREAMBLE_LANE4_END_C = 8'b0;

    localparam QW_IDLE_D = {8{I}};
    localparam QW_IDLE_C = 8'hFF;

    localparam XGMII_ERROR_L0_D = E;
    localparam XGMII_ERROR_L0_C = 8'h01;

    localparam XGMII_ERROR_L4_D = E;
    localparam XGMII_ERROR_L4_C = 8'h10;

    localparam CRC802_3_PRESET = 32'hFFFFFFFF;

    ////////////////////////////////////////////////
    // sof_lane0
    ////////////////////////////////////////////////
    function sof_lane0 (
        input        [63:0]      xgmii_d,
        input        [7:0]       xgmii_c
        );
    begin
        if ((xgmii_d[7:0] == S) && xgmii_c[0])
            sof_lane0 = 1'b1;
        else
            sof_lane0 = 1'b0;
    end
    endfunction // sof_lane0

    ////////////////////////////////////////////////
    // sof_lane0_32
    ////////////////////////////////////////////////
    function sof_lane0_32 (
        input        [31:0]      xgmii_d,
        input        [3:0]       xgmii_c
        );
    begin
        if ((xgmii_d[7:0] == S) && xgmii_c[0])
            sof_lane0_32 = 1'b1;
        else
            sof_lane0_32 = 1'b0;
    end
    endfunction // sof_lane0_32

    ////////////////////////////////////////////////
    // sof_lane4
    ////////////////////////////////////////////////
    function sof_lane4 (
        input        [63:0]      xgmii_d,
        input        [7:0]       xgmii_c
        );
    begin
        if ((xgmii_d[39:32] == S) && xgmii_c[4])
            sof_lane4 = 1'b1;
        else
            sof_lane4 = 1'b0;
    end
    endfunction // sof_lane4

    ////////////////////////////////////////////////
    // crc_rev
    ////////////////////////////////////////////////
    function [31:0] crc_rev (
        input        [31:0]      crc
        );
    integer i;
    reg          [31:0]      o;
    begin
        for (i = 0; i < 32; i = i + 1) begin
            o[i] = crc[31-i];
        end
        crc_rev = o;
    end
    endfunction // crc_rev

    ////////////////////////////////////////////////
    // byte_rev
    ////////////////////////////////////////////////
    function [7:0] byte_rev (
        input        [7:0]       b
        );
    integer i;
    reg          [7:0]       o;
    begin
        for (i = 0; i < 8; i = i + 1) begin
            o[i] = b[7-i];
        end
        byte_rev = o;
    end
    endfunction // byte_rev

    ////////////////////////////////////////////////
    // is_tchar
    ////////////////////////////////////////////////
    function is_tchar (
        input        [7:0]       byte
        );
    begin
        if (byte == T)
            is_tchar = 1'b1;
        else
            is_tchar = 1'b0;
    end
    endfunction // is_tchar

    ////////////////////////////////////////////////
    // crc8B
    ////////////////////////////////////////////////
    function [31:0] crc8B (
        input        [31:0]      c,
        input        [63:0]      d
        );
    reg          [31:0]      o;
    begin
o[0] = d[15] ^ c[12] ^ d[63] ^ d[47] ^ d[39] ^ d[5] ^ d[32] ^ c[28] ^ d[16] ^ c[21] ^ c[13] ^ c[0] ^ d[33] ^ c[29] ^ c[22] ^ d[10] ^ d[57] ^ d[34] ^ d[0] ^ d[26] ^ c[31] ^ d[18] ^ c[23] ^ c[15] ^ d[51] ^ c[2] ^ d[8] ^ d[35] ^ d[19] ^ c[16] ^ d[9] ^ d[2] ^ d[13] ^ d[53] ^ d[37] ^ d[3] ^ d[29] ^ c[26] ^ c[18] ^ d[54] ^ c[5] ^ d[38] ^ d[31] ;
o[1] = c[27] ^ c[19] ^ c[12] ^ d[63] ^ c[6] ^ d[47] ^ d[39] ^ d[5] ^ c[28] ^ d[16] ^ c[21] ^ d[56] ^ d[25] ^ c[30] ^ d[17] ^ d[10] ^ c[14] ^ d[57] ^ d[50] ^ c[1] ^ d[7] ^ d[0] ^ d[26] ^ c[31] ^ c[15] ^ d[51] ^ c[2] ^ d[35] ^ d[1] ^ d[19] ^ d[12] ^ c[24] ^ d[52] ^ c[3] ^ d[36] ^ d[28] ^ d[13] ^ c[17] ^ d[3] ^ d[30] ^ d[29] ^ c[26] ^ d[14] ^ c[18] ^ d[62] ^ d[54] ^ c[5] ^ d[46] ^ d[4] ;
o[2] = c[27] ^ c[19] ^ c[20] ^ c[12] ^ d[63] ^ d[55] ^ c[6] ^ d[47] ^ d[39] ^ d[5] ^ d[32] ^ d[24] ^ c[21] ^ d[56] ^ c[7] ^ c[0] ^ d[33] ^ d[6] ^ d[25] ^ d[10] ^ d[57] ^ d[50] ^ d[49] ^ d[26] ^ d[11] ^ c[23] ^ d[8] ^ d[27] ^ d[19] ^ d[12] ^ c[3] ^ d[28] ^ c[25] ^ d[61] ^ d[45] ^ c[4] ^ d[37] ^ c[26] ^ d[62] ^ d[54] ^ c[5] ^ d[46] ^ d[4] ^ d[31] ;
o[3] = d[23] ^ c[27] ^ c[20] ^ d[55] ^ c[6] ^ d[32] ^ d[5] ^ d[24] ^ c[28] ^ c[21] ^ c[13] ^ d[56] ^ c[7] ^ d[48] ^ c[0] ^ d[25] ^ d[10] ^ c[22] ^ c[8] ^ d[49] ^ c[1] ^ d[7] ^ d[26] ^ d[18] ^ d[11] ^ d[27] ^ c[24] ^ d[60] ^ d[44] ^ d[9] ^ d[36] ^ d[61] ^ d[53] ^ c[4] ^ d[45] ^ d[3] ^ d[30] ^ c[26] ^ d[62] ^ d[54] ^ c[5] ^ d[46] ^ d[38] ^ d[4] ^ d[31] ;
o[4] = d[23] ^ d[15] ^ c[27] ^ c[12] ^ d[63] ^ d[55] ^ c[6] ^ d[39] ^ d[5] ^ d[32] ^ d[24] ^ d[16] ^ c[13] ^ c[7] ^ d[48] ^ d[33] ^ d[6] ^ d[25] ^ d[17] ^ c[14] ^ d[57] ^ c[8] ^ c[1] ^ d[34] ^ d[0] ^ c[31] ^ d[18] ^ c[15] ^ d[51] ^ c[9] ^ d[43] ^ d[19] ^ c[16] ^ d[60] ^ d[59] ^ d[52] ^ d[44] ^ c[25] ^ d[13] ^ d[61] ^ d[45] ^ d[30] ^ d[22] ^ c[26] ^ c[18] ^ d[38] ^ d[4] ;
o[5] = d[23] ^ c[27] ^ c[19] ^ c[12] ^ d[63] ^ d[39] ^ d[24] ^ c[21] ^ d[56] ^ c[7] ^ c[29] ^ d[17] ^ c[22] ^ d[10] ^ c[14] ^ d[57] ^ c[8] ^ d[50] ^ d[42] ^ d[34] ^ d[0] ^ d[26] ^ c[31] ^ c[23] ^ d[58] ^ c[9] ^ d[43] ^ d[8] ^ d[35] ^ d[19] ^ d[12] ^ d[60] ^ d[59] ^ d[44] ^ d[9] ^ d[2] ^ d[21] ^ d[13] ^ c[17] ^ c[10] ^ d[53] ^ d[22] ^ d[14] ^ c[18] ^ d[62] ^ c[5] ^ d[4] ;
o[6] = d[23] ^ c[20] ^ c[19] ^ d[55] ^ c[6] ^ d[16] ^ c[28] ^ c[13] ^ d[56] ^ d[41] ^ d[33] ^ d[25] ^ c[30] ^ c[22] ^ d[57] ^ c[8] ^ d[49] ^ d[42] ^ d[7] ^ d[34] ^ d[18] ^ c[23] ^ d[11] ^ c[15] ^ d[58] ^ c[9] ^ d[43] ^ d[8] ^ d[1] ^ d[20] ^ c[24] ^ d[12] ^ d[59] ^ d[52] ^ d[9] ^ d[21] ^ d[13] ^ c[10] ^ d[61] ^ d[3] ^ d[22] ^ c[18] ^ c[11] ^ d[62] ^ d[38] ;
o[7] = c[19] ^ c[20] ^ d[63] ^ d[55] ^ d[47] ^ d[39] ^ d[40] ^ d[5] ^ d[24] ^ c[28] ^ d[16] ^ c[13] ^ d[56] ^ c[7] ^ d[48] ^ d[41] ^ c[0] ^ d[6] ^ d[17] ^ c[22] ^ c[14] ^ d[42] ^ d[7] ^ d[34] ^ d[26] ^ d[18] ^ d[11] ^ c[15] ^ d[58] ^ c[9] ^ c[2] ^ d[35] ^ d[20] ^ d[12] ^ c[24] ^ d[60] ^ d[9] ^ d[21] ^ c[25] ^ d[13] ^ c[10] ^ d[61] ^ d[53] ^ d[3] ^ d[29] ^ d[22] ^ c[26] ^ c[18] ^ c[11] ^ c[5] ^ d[38] ^ d[31] ;
o[8] = d[23] ^ c[27] ^ c[19] ^ c[20] ^ d[63] ^ d[55] ^ c[6] ^ d[40] ^ d[32] ^ c[28] ^ c[13] ^ d[41] ^ c[0] ^ d[6] ^ d[25] ^ d[17] ^ c[22] ^ c[14] ^ c[8] ^ c[1] ^ d[0] ^ d[26] ^ c[31] ^ d[18] ^ d[11] ^ d[51] ^ c[2] ^ d[35] ^ d[20] ^ d[12] ^ d[60] ^ d[59] ^ d[52] ^ c[3] ^ d[9] ^ d[28] ^ d[21] ^ c[25] ^ d[13] ^ c[10] ^ d[53] ^ d[3] ^ d[30] ^ d[29] ^ c[18] ^ c[11] ^ d[62] ^ c[5] ^ d[46] ^ d[4] ^ d[31] ;
o[9] = c[20] ^ c[19] ^ c[12] ^ c[6] ^ d[40] ^ d[39] ^ d[5] ^ d[24] ^ d[16] ^ c[28] ^ c[21] ^ c[7] ^ c[0] ^ d[25] ^ c[29] ^ d[17] ^ d[10] ^ c[14] ^ d[50] ^ c[1] ^ d[34] ^ c[23] ^ d[11] ^ c[15] ^ d[58] ^ c[9] ^ d[51] ^ c[2] ^ d[8] ^ d[27] ^ d[20] ^ d[19] ^ d[12] ^ d[59] ^ d[52] ^ c[3] ^ d[2] ^ d[28] ^ d[61] ^ c[4] ^ d[45] ^ d[3] ^ d[29] ^ d[30] ^ d[22] ^ c[26] ^ c[11] ^ d[62] ^ d[54] ^ d[31] ;
o[10] = d[23] ^ c[27] ^ c[20] ^ d[63] ^ d[47] ^ d[5] ^ d[32] ^ d[24] ^ c[28] ^ c[7] ^ c[0] ^ c[30] ^ c[8] ^ d[49] ^ d[50] ^ c[1] ^ d[7] ^ d[34] ^ d[0] ^ c[31] ^ d[11] ^ c[23] ^ d[58] ^ d[8] ^ d[35] ^ d[27] ^ d[1] ^ c[24] ^ d[60] ^ c[3] ^ d[44] ^ d[28] ^ d[21] ^ d[13] ^ c[10] ^ d[61] ^ c[4] ^ d[37] ^ d[3] ^ d[30] ^ c[26] ^ c[18] ^ d[54] ^ d[4] ^ d[31] ;
o[11] = d[23] ^ d[15] ^ c[27] ^ c[19] ^ c[12] ^ d[63] ^ d[47] ^ d[39] ^ d[5] ^ d[32] ^ d[16] ^ c[13] ^ d[48] ^ d[6] ^ c[22] ^ c[8] ^ d[49] ^ c[1] ^ d[7] ^ d[18] ^ c[23] ^ c[15] ^ d[51] ^ c[9] ^ d[43] ^ d[8] ^ d[35] ^ d[27] ^ d[20] ^ d[19] ^ d[12] ^ c[24] ^ c[16] ^ d[60] ^ d[59] ^ d[9] ^ d[36] ^ c[25] ^ d[13] ^ c[4] ^ d[37] ^ d[30] ^ d[22] ^ c[26] ^ c[18] ^ c[11] ^ d[62] ^ d[54] ^ d[46] ^ d[38] ^ d[4] ;
o[12] = c[27] ^ c[19] ^ c[20] ^ d[63] ^ d[39] ^ d[32] ^ d[16] ^ c[21] ^ d[48] ^ d[33] ^ d[6] ^ c[29] ^ d[17] ^ c[22] ^ d[10] ^ c[14] ^ d[57] ^ d[50] ^ d[42] ^ d[7] ^ d[0] ^ c[31] ^ d[11] ^ c[15] ^ d[58] ^ d[51] ^ c[9] ^ d[12] ^ c[24] ^ d[59] ^ d[9] ^ d[36] ^ d[2] ^ d[21] ^ c[25] ^ d[13] ^ c[17] ^ c[10] ^ d[61] ^ d[45] ^ d[22] ^ d[14] ^ c[18] ^ d[62] ^ d[54] ^ d[46] ^ d[4] ;
o[13] = d[15] ^ c[20] ^ c[19] ^ d[47] ^ d[32] ^ d[5] ^ d[16] ^ c[28] ^ c[21] ^ d[56] ^ d[41] ^ c[0] ^ d[6] ^ c[30] ^ d[10] ^ c[22] ^ d[57] ^ d[50] ^ d[49] ^ c[23] ^ d[11] ^ c[15] ^ d[58] ^ d[8] ^ d[35] ^ d[1] ^ d[20] ^ d[12] ^ c[16] ^ d[60] ^ d[44] ^ d[9] ^ d[21] ^ c[25] ^ d[13] ^ c[10] ^ d[61] ^ d[53] ^ d[45] ^ d[3] ^ c[26] ^ c[18] ^ c[11] ^ d[62] ^ d[38] ^ d[31] ;
o[14] = c[27] ^ d[15] ^ c[19] ^ c[20] ^ c[12] ^ d[55] ^ d[40] ^ d[5] ^ c[21] ^ d[56] ^ d[48] ^ c[0] ^ c[29] ^ d[10] ^ c[22] ^ d[57] ^ d[49] ^ c[1] ^ d[7] ^ d[34] ^ d[0] ^ c[31] ^ d[11] ^ c[23] ^ d[43] ^ d[8] ^ d[19] ^ d[20] ^ c[24] ^ d[12] ^ c[16] ^ d[60] ^ d[59] ^ d[52] ^ d[44] ^ d[9] ^ d[2] ^ c[17] ^ d[61] ^ d[37] ^ d[30] ^ c[26] ^ d[14] ^ c[11] ^ d[46] ^ d[31] ^ d[4] ;
o[15] = c[27] ^ c[20] ^ c[12] ^ d[55] ^ d[47] ^ d[39] ^ c[28] ^ c[21] ^ c[13] ^ d[56] ^ d[48] ^ d[6] ^ d[33] ^ c[30] ^ c[22] ^ d[10] ^ d[42] ^ c[1] ^ d[7] ^ d[18] ^ c[23] ^ d[11] ^ d[58] ^ d[51] ^ c[2] ^ d[43] ^ d[8] ^ d[1] ^ d[19] ^ c[24] ^ d[60] ^ d[59] ^ d[36] ^ d[9] ^ c[25] ^ d[13] ^ c[17] ^ d[45] ^ d[30] ^ d[3] ^ d[29] ^ d[14] ^ c[18] ^ d[54] ^ d[4] ;
o[16] = d[15] ^ c[19] ^ c[12] ^ d[63] ^ d[55] ^ d[39] ^ d[16] ^ d[41] ^ c[0] ^ d[33] ^ d[6] ^ d[17] ^ c[14] ^ d[50] ^ d[42] ^ d[7] ^ d[34] ^ d[26] ^ c[15] ^ d[58] ^ d[51] ^ d[19] ^ d[12] ^ c[24] ^ c[16] ^ d[59] ^ c[3] ^ d[44] ^ d[28] ^ c[25] ^ d[37] ^ c[5] ^ d[46] ^ d[31] ;
o[17] = d[15] ^ c[20] ^ c[6] ^ d[40] ^ d[32] ^ d[5] ^ d[16] ^ c[13] ^ d[41] ^ d[6] ^ d[33] ^ d[25] ^ d[57] ^ d[50] ^ d[49] ^ c[1] ^ d[18] ^ d[11] ^ c[15] ^ d[58] ^ d[43] ^ d[27] ^ c[16] ^ d[36] ^ c[25] ^ c[17] ^ c[4] ^ d[45] ^ d[30] ^ d[14] ^ c[26] ^ d[62] ^ d[54] ^ d[38] ;
o[18] = c[27] ^ d[15] ^ d[40] ^ d[39] ^ d[5] ^ d[32] ^ d[24] ^ c[21] ^ d[56] ^ c[7] ^ d[48] ^ c[0] ^ d[17] ^ d[10] ^ c[14] ^ d[57] ^ d[49] ^ d[42] ^ d[26] ^ c[2] ^ d[35] ^ c[16] ^ d[44] ^ d[13] ^ c[17] ^ d[61] ^ d[53] ^ d[37] ^ d[29] ^ c[26] ^ d[14] ^ c[18] ^ c[5] ^ d[31] ^ d[4] ;
o[19] = d[23] ^ c[27] ^ c[19] ^ d[55] ^ c[6] ^ d[47] ^ d[39] ^ c[28] ^ d[16] ^ d[56] ^ d[48] ^ d[41] ^ c[0] ^ d[25] ^ c[22] ^ c[8] ^ c[1] ^ d[34] ^ c[15] ^ d[43] ^ d[12] ^ d[60] ^ d[52] ^ c[3] ^ d[36] ^ d[9] ^ d[28] ^ d[13] ^ c[17] ^ d[30] ^ d[3] ^ d[14] ^ c[18] ^ d[38] ^ d[4] ^ d[31] ;
o[20] = d[15] ^ c[20] ^ c[19] ^ d[55] ^ d[47] ^ d[40] ^ d[24] ^ c[28] ^ c[7] ^ d[33] ^ c[29] ^ c[1] ^ d[42] ^ d[11] ^ c[23] ^ c[9] ^ d[51] ^ c[2] ^ d[35] ^ d[8] ^ d[27] ^ d[12] ^ c[16] ^ d[59] ^ d[2] ^ d[13] ^ c[4] ^ d[37] ^ d[29] ^ d[3] ^ d[30] ^ d[22] ^ c[18] ^ d[54] ^ d[46] ^ d[38] ;
o[21] = d[23] ^ c[19] ^ c[20] ^ d[39] ^ d[32] ^ c[21] ^ d[41] ^ c[30] ^ c[29] ^ d[10] ^ c[8] ^ d[50] ^ d[34] ^ d[7] ^ d[26] ^ d[11] ^ d[58] ^ c[2] ^ d[1] ^ c[24] ^ d[12] ^ c[3] ^ d[36] ^ d[28] ^ d[2] ^ d[21] ^ c[17] ^ c[10] ^ d[53] ^ d[45] ^ d[37] ^ d[29] ^ d[14] ^ d[54] ^ d[46] ^ c[5] ;
o[22] = d[15] ^ c[20] ^ c[12] ^ d[63] ^ c[6] ^ d[47] ^ d[39] ^ d[40] ^ d[5] ^ d[32] ^ c[28] ^ d[16] ^ c[13] ^ d[6] ^ d[25] ^ c[29] ^ c[30] ^ d[49] ^ d[34] ^ d[26] ^ d[18] ^ d[11] ^ c[23] ^ c[15] ^ d[51] ^ c[9] ^ c[2] ^ d[8] ^ d[27] ^ d[1] ^ d[20] ^ d[19] ^ c[16] ^ d[52] ^ c[3] ^ d[44] ^ d[36] ^ d[2] ^ d[28] ^ c[25] ^ d[45] ^ c[4] ^ d[37] ^ d[3] ^ d[29] ^ d[22] ^ c[26] ^ c[11] ^ d[54] ^ c[5] ;
o[23] = c[27] ^ d[63] ^ c[6] ^ d[47] ^ d[32] ^ d[24] ^ c[28] ^ d[16] ^ c[7] ^ d[48] ^ d[25] ^ c[30] ^ d[17] ^ c[22] ^ c[14] ^ d[57] ^ d[50] ^ d[7] ^ d[34] ^ c[23] ^ c[15] ^ c[2] ^ d[43] ^ d[8] ^ d[27] ^ d[1] ^ c[24] ^ c[3] ^ d[44] ^ d[9] ^ d[36] ^ d[28] ^ d[21] ^ d[13] ^ c[17] ^ c[10] ^ c[4] ^ d[37] ^ d[3] ^ d[29] ^ d[14] ^ c[18] ^ d[62] ^ d[54] ^ d[46] ^ d[4] ;
o[24] = d[23] ^ d[15] ^ c[19] ^ d[47] ^ d[24] ^ d[16] ^ c[28] ^ d[56] ^ c[7] ^ c[0] ^ d[6] ^ d[33] ^ c[29] ^ c[8] ^ d[49] ^ d[42] ^ d[7] ^ d[26] ^ d[0] ^ c[31] ^ c[23] ^ c[15] ^ d[43] ^ d[8] ^ d[35] ^ d[27] ^ d[20] ^ c[24] ^ d[12] ^ c[16] ^ c[3] ^ d[36] ^ d[2] ^ d[28] ^ c[25] ^ d[13] ^ d[61] ^ d[53] ^ c[4] ^ d[45] ^ d[3] ^ c[18] ^ c[11] ^ d[62] ^ c[5] ^ d[46] ^ d[31] ;
o[25] = d[23] ^ d[15] ^ c[19] ^ c[20] ^ c[12] ^ d[55] ^ c[6] ^ d[5] ^ d[32] ^ d[48] ^ d[41] ^ d[6] ^ d[25] ^ c[30] ^ c[29] ^ c[8] ^ c[1] ^ d[42] ^ d[7] ^ d[34] ^ d[26] ^ d[11] ^ c[9] ^ d[35] ^ d[1] ^ d[27] ^ d[19] ^ c[24] ^ d[12] ^ c[16] ^ d[60] ^ d[52] ^ d[44] ^ d[2] ^ c[25] ^ c[17] ^ d[61] ^ c[4] ^ d[45] ^ d[30] ^ d[22] ^ c[26] ^ d[14] ^ d[46] ^ c[5] ;
o[26] = d[15] ^ c[27] ^ c[20] ^ c[12] ^ d[63] ^ c[6] ^ d[39] ^ d[40] ^ d[32] ^ d[24] ^ c[28] ^ d[16] ^ c[7] ^ d[41] ^ d[6] ^ d[25] ^ c[29] ^ c[30] ^ c[22] ^ d[57] ^ d[11] ^ c[23] ^ c[15] ^ c[9] ^ d[43] ^ d[8] ^ d[35] ^ d[1] ^ d[19] ^ c[16] ^ d[60] ^ d[59] ^ d[44] ^ d[9] ^ d[2] ^ d[21] ^ c[25] ^ c[17] ^ c[10] ^ d[53] ^ d[45] ^ d[37] ^ d[3] ^ d[22] ^ d[14] ^ d[38] ^ d[4] ;
o[27] = d[23] ^ d[15] ^ d[40] ^ d[39] ^ d[5] ^ d[24] ^ c[28] ^ c[21] ^ c[13] ^ d[56] ^ c[7] ^ c[0] ^ c[29] ^ c[30] ^ d[10] ^ c[8] ^ d[42] ^ d[7] ^ d[34] ^ d[0] ^ c[31] ^ d[18] ^ c[23] ^ d[58] ^ d[43] ^ d[8] ^ d[1] ^ d[20] ^ c[24] ^ c[16] ^ d[59] ^ d[52] ^ d[44] ^ d[36] ^ d[2] ^ d[21] ^ d[13] ^ c[17] ^ c[10] ^ d[37] ^ d[3] ^ d[14] ^ c[26] ^ c[18] ^ c[11] ^ d[62] ^ d[38] ^ d[31] ;
o[28] = d[23] ^ c[27] ^ c[19] ^ c[12] ^ d[55] ^ d[39] ^ d[41] ^ d[6] ^ d[33] ^ c[30] ^ c[29] ^ d[17] ^ c[22] ^ c[14] ^ d[57] ^ c[8] ^ c[1] ^ d[42] ^ d[7] ^ d[0] ^ c[31] ^ d[58] ^ c[9] ^ d[51] ^ d[43] ^ d[35] ^ d[1] ^ d[19] ^ d[20] ^ c[24] ^ d[12] ^ d[9] ^ d[36] ^ d[2] ^ d[13] ^ c[25] ^ c[17] ^ d[61] ^ d[37] ^ d[30] ^ d[22] ^ d[14] ^ c[18] ^ c[11] ^ d[38] ^ d[4] ;
o[29] = c[19] ^ c[20] ^ c[12] ^ d[40] ^ d[5] ^ d[32] ^ c[28] ^ d[16] ^ c[13] ^ d[56] ^ d[41] ^ d[6] ^ c[30] ^ d[57] ^ d[50] ^ d[42] ^ d[34] ^ d[0] ^ d[18] ^ c[31] ^ c[23] ^ d[11] ^ c[15] ^ c[9] ^ c[2] ^ d[8] ^ d[35] ^ d[1] ^ d[19] ^ d[12] ^ d[60] ^ d[36] ^ d[21] ^ c[25] ^ d[13] ^ c[10] ^ d[37] ^ d[3] ^ d[29] ^ d[22] ^ c[26] ^ c[18] ^ d[54] ^ d[38] ;
o[30] = c[27] ^ d[15] ^ c[20] ^ c[19] ^ d[55] ^ d[40] ^ d[39] ^ d[5] ^ c[21] ^ c[13] ^ d[56] ^ d[41] ^ c[0] ^ d[33] ^ d[17] ^ c[29] ^ d[10] ^ c[14] ^ d[49] ^ d[7] ^ d[34] ^ d[0] ^ c[31] ^ d[18] ^ d[11] ^ d[35] ^ d[20] ^ c[24] ^ d[12] ^ c[16] ^ d[59] ^ c[3] ^ d[36] ^ d[2] ^ d[28] ^ d[21] ^ c[10] ^ d[53] ^ d[37] ^ c[26] ^ c[11] ^ d[4] ^ d[31] ;
o[31] = c[27] ^ c[20] ^ c[12] ^ d[55] ^ d[40] ^ d[39] ^ d[32] ^ d[16] ^ c[28] ^ c[21] ^ d[48] ^ d[6] ^ d[33] ^ c[30] ^ d[17] ^ d[10] ^ c[22] ^ c[14] ^ c[1] ^ d[34] ^ d[11] ^ c[15] ^ d[58] ^ d[35] ^ d[1] ^ d[27] ^ d[19] ^ d[20] ^ d[52] ^ d[9] ^ d[36] ^ c[25] ^ c[17] ^ c[4] ^ d[3] ^ d[30] ^ d[14] ^ c[11] ^ d[54] ^ d[38] ^ d[4] ;
        crc8B = o;
    end
    endfunction // crc8B

    ////////////////////////////////////////////////
    // crc7B
    ////////////////////////////////////////////////
    function [31:0] crc7B (
        input        [31:0]      c,
        input        [55:0]      d
        );
    reg          [31:0]      o;
    begin
o[0] = d[23] ^ c[20] ^ d[55] ^ c[6] ^ d[39] ^ d[5] ^ d[24] ^ c[21] ^ c[13] ^ c[7] ^ c[0] ^ d[25] ^ c[30] ^ c[29] ^ d[10] ^ d[49] ^ c[8] ^ c[1] ^ d[7] ^ d[0] ^ d[26] ^ c[31] ^ d[18] ^ d[11] ^ c[23] ^ d[43] ^ c[2] ^ d[8] ^ d[1] ^ d[27] ^ c[24] ^ d[2] ^ d[21] ^ c[10] ^ c[4] ^ d[45] ^ d[30] ^ d[29] ^ c[26] ^ d[46] ^ c[5] ^ d[31] ;
o[1] = c[27] ^ c[20] ^ d[55] ^ d[39] ^ d[5] ^ c[13] ^ d[48] ^ c[0] ^ d[6] ^ c[29] ^ d[17] ^ c[22] ^ c[14] ^ d[49] ^ d[42] ^ d[18] ^ d[11] ^ c[23] ^ c[9] ^ d[43] ^ d[8] ^ d[27] ^ d[20] ^ c[3] ^ d[44] ^ d[9] ^ d[2] ^ d[28] ^ d[21] ^ c[25] ^ c[10] ^ c[4] ^ d[22] ^ c[26] ^ c[11] ^ d[54] ^ d[46] ^ d[38] ^ d[31] ^ d[4] ;
o[2] = d[23] ^ c[27] ^ c[20] ^ c[12] ^ d[55] ^ c[6] ^ d[47] ^ d[39] ^ d[24] ^ c[28] ^ d[16] ^ c[13] ^ c[7] ^ d[48] ^ c[0] ^ d[41] ^ d[25] ^ c[29] ^ d[17] ^ c[14] ^ d[49] ^ c[8] ^ d[42] ^ d[0] ^ c[31] ^ d[18] ^ d[11] ^ c[15] ^ c[2] ^ d[19] ^ d[20] ^ d[2] ^ d[53] ^ d[37] ^ d[3] ^ d[29] ^ c[11] ^ d[54] ^ d[46] ^ d[38] ^ d[31] ^ d[4] ;
o[3] = d[23] ^ d[15] ^ c[12] ^ d[47] ^ d[40] ^ d[24] ^ c[28] ^ d[16] ^ c[21] ^ c[13] ^ d[48] ^ c[7] ^ d[41] ^ c[29] ^ c[30] ^ d[17] ^ d[10] ^ c[14] ^ c[8] ^ c[1] ^ d[18] ^ c[15] ^ c[9] ^ d[1] ^ d[19] ^ c[16] ^ d[52] ^ c[3] ^ d[36] ^ d[2] ^ d[28] ^ d[53] ^ d[45] ^ d[37] ^ d[30] ^ d[3] ^ d[22] ^ d[54] ^ d[46] ^ d[38] ;
o[4] = d[15] ^ c[20] ^ d[55] ^ c[6] ^ d[47] ^ d[40] ^ d[5] ^ d[24] ^ d[16] ^ c[21] ^ c[7] ^ c[0] ^ d[25] ^ d[17] ^ d[10] ^ c[22] ^ c[14] ^ d[49] ^ c[1] ^ d[7] ^ d[26] ^ d[11] ^ c[23] ^ c[15] ^ c[9] ^ d[51] ^ d[43] ^ d[8] ^ d[35] ^ c[24] ^ c[16] ^ d[52] ^ d[44] ^ d[9] ^ d[36] ^ c[17] ^ d[53] ^ d[37] ^ d[30] ^ d[22] ^ c[26] ^ d[14] ^ c[5] ^ d[31] ;
o[5] = c[27] ^ d[15] ^ c[20] ^ d[55] ^ d[5] ^ d[16] ^ c[13] ^ d[48] ^ c[0] ^ d[6] ^ c[30] ^ c[29] ^ c[22] ^ d[49] ^ d[50] ^ d[42] ^ d[34] ^ d[0] ^ d[26] ^ c[31] ^ d[18] ^ d[11] ^ c[15] ^ d[51] ^ d[35] ^ d[1] ^ d[27] ^ c[16] ^ d[52] ^ d[9] ^ d[36] ^ d[2] ^ d[13] ^ c[25] ^ c[17] ^ c[4] ^ d[45] ^ c[26] ^ d[14] ^ c[18] ^ d[54] ^ c[5] ^ d[31] ^ d[4] ;
o[6] = d[15] ^ c[27] ^ c[19] ^ c[6] ^ d[47] ^ d[5] ^ c[28] ^ c[21] ^ d[48] ^ d[41] ^ d[33] ^ d[25] ^ c[30] ^ d[17] ^ d[10] ^ c[14] ^ d[50] ^ d[49] ^ c[1] ^ d[34] ^ d[0] ^ d[26] ^ c[31] ^ c[23] ^ d[51] ^ d[8] ^ d[35] ^ d[1] ^ d[12] ^ c[16] ^ d[44] ^ d[13] ^ c[17] ^ d[53] ^ d[30] ^ d[3] ^ c[26] ^ d[14] ^ c[18] ^ d[54] ^ c[5] ^ d[4] ;
o[7] = d[23] ^ c[27] ^ c[19] ^ d[55] ^ d[47] ^ d[40] ^ d[39] ^ d[5] ^ d[32] ^ c[28] ^ d[16] ^ c[21] ^ c[13] ^ d[48] ^ c[0] ^ d[33] ^ c[30] ^ d[10] ^ c[22] ^ c[8] ^ d[50] ^ c[1] ^ d[34] ^ d[26] ^ d[18] ^ c[23] ^ c[15] ^ d[8] ^ d[1] ^ d[27] ^ d[12] ^ d[52] ^ d[9] ^ d[21] ^ d[13] ^ c[17] ^ c[10] ^ d[53] ^ c[4] ^ d[45] ^ d[3] ^ d[30] ^ c[26] ^ d[14] ^ c[18] ^ c[5] ^ d[31] ^ d[4] ;
o[8] = d[23] ^ c[27] ^ d[15] ^ c[19] ^ d[55] ^ d[47] ^ d[5] ^ d[32] ^ d[24] ^ c[28] ^ c[21] ^ c[13] ^ c[7] ^ d[33] ^ c[30] ^ d[17] ^ d[10] ^ c[22] ^ c[14] ^ c[8] ^ d[18] ^ c[9] ^ d[51] ^ d[43] ^ d[1] ^ d[27] ^ d[20] ^ d[12] ^ c[16] ^ d[52] ^ d[44] ^ d[9] ^ d[21] ^ d[13] ^ c[10] ^ c[4] ^ d[45] ^ d[3] ^ d[22] ^ c[26] ^ c[18] ^ c[11] ^ d[54] ^ d[38] ^ d[4] ;
o[9] = d[23] ^ c[27] ^ c[19] ^ c[20] ^ c[12] ^ d[32] ^ c[28] ^ d[16] ^ c[0] ^ c[29] ^ d[17] ^ c[22] ^ c[14] ^ c[8] ^ d[50] ^ d[42] ^ d[0] ^ d[26] ^ c[31] ^ c[23] ^ d[11] ^ c[15] ^ c[9] ^ d[51] ^ d[43] ^ d[8] ^ d[20] ^ d[19] ^ d[12] ^ d[44] ^ d[9] ^ d[2] ^ d[21] ^ c[17] ^ c[10] ^ d[53] ^ d[37] ^ d[3] ^ d[22] ^ d[14] ^ c[11] ^ d[54] ^ c[5] ^ d[46] ^ d[4] ^ d[31] ;
o[10] = d[23] ^ d[15] ^ c[12] ^ d[55] ^ d[39] ^ d[5] ^ d[24] ^ c[28] ^ d[16] ^ c[7] ^ d[41] ^ c[8] ^ d[50] ^ d[42] ^ d[0] ^ d[26] ^ c[31] ^ c[15] ^ c[9] ^ c[2] ^ d[27] ^ d[19] ^ d[20] ^ c[16] ^ d[52] ^ d[36] ^ d[13] ^ d[53] ^ c[4] ^ d[3] ^ d[29] ^ d[22] ^ c[26] ^ c[18] ^ c[11] ^ d[46] ^ c[5] ;
o[11] = c[27] ^ d[15] ^ c[19] ^ c[20] ^ c[12] ^ d[55] ^ d[40] ^ d[39] ^ d[5] ^ d[24] ^ c[21] ^ c[7] ^ c[0] ^ d[41] ^ c[30] ^ d[10] ^ c[1] ^ d[7] ^ d[0] ^ c[31] ^ d[11] ^ c[23] ^ c[9] ^ d[51] ^ d[43] ^ c[2] ^ d[8] ^ d[35] ^ d[1] ^ d[27] ^ d[19] ^ c[24] ^ d[12] ^ c[16] ^ d[52] ^ c[3] ^ d[28] ^ c[17] ^ c[4] ^ d[30] ^ d[29] ^ d[22] ^ c[26] ^ d[14] ^ d[54] ^ d[46] ^ d[38] ^ d[31] ^ d[4] ;
o[12] = c[27] ^ d[55] ^ c[6] ^ d[40] ^ d[5] ^ d[24] ^ c[28] ^ c[7] ^ c[0] ^ d[6] ^ d[25] ^ c[30] ^ c[29] ^ c[22] ^ d[49] ^ d[50] ^ d[42] ^ d[34] ^ c[23] ^ d[51] ^ d[43] ^ d[8] ^ d[1] ^ c[3] ^ d[9] ^ d[2] ^ d[28] ^ d[13] ^ c[25] ^ c[17] ^ d[53] ^ d[37] ^ d[3] ^ c[26] ^ d[14] ^ c[18] ^ d[54] ^ d[46] ^ d[38] ^ d[31] ^ d[4] ;
o[13] = d[23] ^ c[27] ^ c[19] ^ d[39] ^ d[5] ^ d[24] ^ c[28] ^ d[48] ^ c[7] ^ d[41] ^ d[33] ^ c[29] ^ c[30] ^ c[8] ^ d[50] ^ d[49] ^ d[42] ^ c[1] ^ d[7] ^ d[0] ^ c[31] ^ c[23] ^ d[8] ^ d[1] ^ d[27] ^ d[12] ^ c[24] ^ d[52] ^ d[36] ^ d[2] ^ d[13] ^ d[53] ^ c[4] ^ d[45] ^ d[37] ^ d[30] ^ d[3] ^ c[26] ^ c[18] ^ d[54] ^ d[4] ;
o[14] = d[23] ^ c[27] ^ c[20] ^ c[19] ^ d[47] ^ d[40] ^ d[32] ^ c[28] ^ d[48] ^ d[41] ^ d[6] ^ c[29] ^ c[30] ^ c[8] ^ d[49] ^ d[7] ^ d[0] ^ d[26] ^ c[31] ^ d[11] ^ c[9] ^ d[51] ^ c[2] ^ d[35] ^ d[1] ^ c[24] ^ d[12] ^ d[52] ^ d[44] ^ d[36] ^ d[2] ^ c[25] ^ d[53] ^ d[29] ^ d[3] ^ d[22] ^ c[5] ^ d[38] ^ d[4] ;
o[15] = c[20] ^ c[6] ^ d[47] ^ d[40] ^ d[39] ^ d[5] ^ c[28] ^ c[21] ^ d[48] ^ c[0] ^ d[6] ^ d[25] ^ c[30] ^ c[29] ^ d[10] ^ d[50] ^ d[34] ^ d[0] ^ c[31] ^ d[11] ^ c[9] ^ d[51] ^ d[43] ^ d[35] ^ d[1] ^ d[52] ^ c[3] ^ d[28] ^ d[2] ^ d[21] ^ c[25] ^ c[10] ^ d[37] ^ d[3] ^ d[22] ^ c[26] ^ d[46] ^ d[31] ;
o[16] = d[23] ^ c[27] ^ c[20] ^ d[55] ^ c[6] ^ d[47] ^ c[13] ^ c[0] ^ d[33] ^ d[25] ^ c[22] ^ c[8] ^ d[50] ^ d[42] ^ d[7] ^ d[34] ^ d[26] ^ d[18] ^ d[11] ^ c[23] ^ d[51] ^ d[43] ^ c[2] ^ d[8] ^ d[20] ^ c[24] ^ d[9] ^ d[36] ^ d[29] ^ c[11] ^ c[5] ^ d[38] ^ d[31] ^ d[4] ;
o[17] = c[12] ^ c[6] ^ d[32] ^ d[24] ^ c[28] ^ c[21] ^ c[7] ^ d[41] ^ d[6] ^ d[33] ^ d[25] ^ d[17] ^ d[10] ^ c[14] ^ d[50] ^ d[49] ^ d[42] ^ c[1] ^ d[7] ^ c[23] ^ c[9] ^ d[8] ^ d[35] ^ d[19] ^ c[24] ^ c[3] ^ d[28] ^ c[25] ^ d[37] ^ d[30] ^ d[3] ^ d[22] ^ d[54] ^ d[46] ;
o[18] = d[23] ^ d[40] ^ d[5] ^ d[32] ^ d[24] ^ d[16] ^ c[13] ^ c[7] ^ d[48] ^ d[41] ^ c[0] ^ d[6] ^ c[29] ^ c[22] ^ c[8] ^ d[49] ^ d[7] ^ d[34] ^ d[18] ^ c[15] ^ c[2] ^ d[27] ^ c[24] ^ d[9] ^ d[36] ^ d[2] ^ d[21] ^ c[25] ^ c[10] ^ d[53] ^ c[4] ^ d[45] ^ d[29] ^ c[26] ^ d[31] ;
o[19] = d[23] ^ c[27] ^ d[15] ^ d[47] ^ d[40] ^ d[39] ^ d[5] ^ d[48] ^ c[0] ^ d[6] ^ d[33] ^ c[30] ^ d[17] ^ c[14] ^ c[8] ^ c[1] ^ d[26] ^ c[23] ^ c[9] ^ d[8] ^ d[35] ^ d[1] ^ d[20] ^ c[16] ^ d[52] ^ c[3] ^ d[44] ^ d[28] ^ c[25] ^ d[30] ^ d[22] ^ c[26] ^ c[11] ^ c[5] ^ d[4] ^ d[31] ;
o[20] = c[27] ^ c[12] ^ c[6] ^ d[47] ^ d[39] ^ d[5] ^ d[32] ^ c[28] ^ d[16] ^ d[25] ^ c[1] ^ d[7] ^ d[34] ^ d[0] ^ c[31] ^ c[15] ^ d[51] ^ c[9] ^ c[2] ^ d[43] ^ d[27] ^ d[19] ^ c[24] ^ d[21] ^ c[17] ^ c[10] ^ c[4] ^ d[3] ^ d[30] ^ d[29] ^ d[22] ^ c[26] ^ d[14] ^ d[46] ^ d[38] ^ d[4] ;
o[21] = c[27] ^ d[15] ^ d[24] ^ c[28] ^ c[13] ^ c[7] ^ c[0] ^ d[6] ^ d[33] ^ c[29] ^ d[50] ^ d[42] ^ d[26] ^ d[18] ^ c[2] ^ d[20] ^ c[16] ^ c[3] ^ d[2] ^ d[28] ^ d[21] ^ c[25] ^ d[13] ^ c[10] ^ d[45] ^ d[37] ^ d[3] ^ d[29] ^ c[18] ^ c[11] ^ c[5] ^ d[46] ^ d[38] ^ d[4] ^ d[31] ;
o[22] = c[19] ^ c[20] ^ c[12] ^ d[55] ^ d[39] ^ d[32] ^ d[24] ^ c[28] ^ c[21] ^ c[13] ^ c[7] ^ c[0] ^ d[41] ^ d[17] ^ d[10] ^ c[14] ^ d[7] ^ d[0] ^ d[26] ^ c[31] ^ d[18] ^ d[11] ^ c[23] ^ d[43] ^ c[2] ^ d[8] ^ d[19] ^ d[20] ^ c[24] ^ d[12] ^ c[3] ^ d[44] ^ d[36] ^ d[28] ^ d[21] ^ c[17] ^ c[10] ^ d[37] ^ d[3] ^ d[29] ^ d[14] ^ c[11] ^ d[46] ^ c[5] ^ d[31] ;
o[23] = c[12] ^ d[55] ^ d[40] ^ d[39] ^ d[5] ^ d[24] ^ d[16] ^ c[7] ^ d[6] ^ c[30] ^ d[17] ^ c[22] ^ c[14] ^ d[49] ^ d[42] ^ d[0] ^ d[26] ^ c[31] ^ c[23] ^ c[15] ^ c[2] ^ d[8] ^ d[35] ^ d[1] ^ d[19] ^ d[20] ^ c[3] ^ d[9] ^ d[36] ^ d[28] ^ d[21] ^ d[13] ^ c[25] ^ c[10] ^ d[29] ^ c[26] ^ c[18] ^ c[11] ^ d[54] ^ d[46] ^ c[5] ^ d[38] ;
o[24] = d[23] ^ d[15] ^ c[27] ^ c[19] ^ c[12] ^ c[6] ^ d[39] ^ d[5] ^ d[16] ^ c[13] ^ d[48] ^ d[41] ^ d[25] ^ c[8] ^ d[7] ^ d[34] ^ d[0] ^ d[18] ^ c[31] ^ c[23] ^ c[15] ^ d[8] ^ d[35] ^ d[27] ^ d[20] ^ d[19] ^ d[12] ^ c[24] ^ c[16] ^ c[3] ^ d[28] ^ d[53] ^ c[4] ^ d[45] ^ d[37] ^ c[26] ^ c[11] ^ d[54] ^ d[38] ^ d[4] ;
o[25] = c[27] ^ d[15] ^ c[20] ^ c[12] ^ d[47] ^ d[40] ^ d[24] ^ c[28] ^ c[13] ^ c[7] ^ d[6] ^ d[33] ^ d[17] ^ c[14] ^ d[7] ^ d[34] ^ d[26] ^ d[18] ^ d[11] ^ c[9] ^ d[27] ^ d[19] ^ c[24] ^ c[16] ^ d[52] ^ d[44] ^ d[36] ^ c[25] ^ c[17] ^ d[53] ^ c[4] ^ d[37] ^ d[3] ^ d[22] ^ d[14] ^ c[5] ^ d[38] ^ d[4] ;
o[26] = c[20] ^ d[55] ^ d[32] ^ d[24] ^ c[28] ^ d[16] ^ c[7] ^ c[0] ^ d[6] ^ d[33] ^ c[30] ^ d[17] ^ c[14] ^ d[49] ^ c[1] ^ d[7] ^ d[0] ^ c[31] ^ d[11] ^ c[23] ^ c[15] ^ d[51] ^ c[2] ^ d[8] ^ d[35] ^ d[1] ^ d[27] ^ c[24] ^ d[52] ^ d[36] ^ d[13] ^ c[25] ^ c[17] ^ c[4] ^ d[45] ^ d[37] ^ d[3] ^ d[30] ^ d[29] ^ d[14] ^ c[18] ^ d[31] ;
o[27] = d[23] ^ d[15] ^ c[19] ^ d[5] ^ d[32] ^ d[16] ^ c[21] ^ d[48] ^ c[0] ^ d[6] ^ c[29] ^ d[10] ^ c[8] ^ d[50] ^ c[1] ^ d[7] ^ d[34] ^ d[0] ^ d[26] ^ c[31] ^ c[15] ^ d[51] ^ c[2] ^ d[35] ^ d[12] ^ c[24] ^ c[16] ^ c[3] ^ d[44] ^ d[36] ^ d[2] ^ d[28] ^ c[25] ^ d[13] ^ d[30] ^ d[29] ^ c[26] ^ c[18] ^ d[54] ^ c[5] ^ d[31] ;
o[28] = c[27] ^ d[15] ^ c[20] ^ c[19] ^ d[47] ^ c[6] ^ d[5] ^ c[0] ^ d[6] ^ d[33] ^ d[25] ^ c[30] ^ c[22] ^ d[50] ^ d[49] ^ c[1] ^ d[34] ^ d[11] ^ c[9] ^ c[2] ^ d[43] ^ d[35] ^ d[1] ^ d[27] ^ d[12] ^ c[16] ^ c[3] ^ d[9] ^ d[28] ^ c[25] ^ c[17] ^ d[53] ^ c[4] ^ d[29] ^ d[30] ^ d[22] ^ c[26] ^ d[14] ^ d[4] ^ d[31] ;
o[29] = c[27] ^ c[20] ^ d[5] ^ d[32] ^ d[24] ^ c[28] ^ c[21] ^ c[7] ^ d[48] ^ d[33] ^ d[10] ^ d[49] ^ c[1] ^ d[42] ^ d[34] ^ d[0] ^ d[26] ^ c[31] ^ c[23] ^ d[11] ^ c[2] ^ d[8] ^ d[27] ^ d[52] ^ c[3] ^ d[28] ^ d[21] ^ d[13] ^ c[17] ^ c[10] ^ c[4] ^ d[3] ^ d[30] ^ d[29] ^ c[26] ^ d[14] ^ c[18] ^ d[46] ^ c[5] ^ d[4] ;
o[30] = d[23] ^ c[27] ^ c[19] ^ c[6] ^ d[47] ^ d[32] ^ c[28] ^ c[21] ^ d[48] ^ d[41] ^ c[0] ^ d[33] ^ d[25] ^ c[29] ^ c[22] ^ d[10] ^ c[8] ^ d[7] ^ d[26] ^ d[51] ^ c[2] ^ d[27] ^ d[20] ^ d[12] ^ c[24] ^ c[3] ^ d[9] ^ d[2] ^ d[28] ^ d[13] ^ d[45] ^ c[4] ^ d[3] ^ d[29] ^ c[18] ^ c[11] ^ c[5] ^ d[4] ^ d[31] ;
o[31] = c[20] ^ c[19] ^ c[12] ^ c[6] ^ d[47] ^ d[40] ^ d[32] ^ d[24] ^ c[28] ^ c[7] ^ c[0] ^ d[6] ^ d[25] ^ c[29] ^ c[30] ^ c[22] ^ d[50] ^ c[1] ^ d[26] ^ c[23] ^ d[11] ^ c[9] ^ d[8] ^ d[1] ^ d[27] ^ d[19] ^ d[12] ^ d[44] ^ c[3] ^ d[9] ^ d[2] ^ d[28] ^ c[25] ^ c[4] ^ d[3] ^ d[30] ^ d[22] ^ c[5] ^ d[46] ^ d[31] ;
        crc7B = o;
    end
    endfunction // crc7B

    ////////////////////////////////////////////////
    // crc6B
    ////////////////////////////////////////////////
    function [31:0] crc6B (
        input        [31:0]      c,
        input        [47:0]      d
        );
    reg          [31:0]      o;
    begin
o[0] = d[41] ^ d[23] ^ c[0] ^ d[15] ^ c[9] ^ c[10] ^ d[35] ^ d[17] ^ c[29] ^ c[12] ^ d[10] ^ c[14] ^ d[19] ^ d[37] ^ d[47] ^ d[3] ^ c[16] ^ d[22] ^ c[8] ^ c[18] ^ c[28] ^ d[16] ^ d[0] ^ c[21] ^ c[31] ^ d[18] ^ c[13] ^ d[2] ^ c[15] ^ d[21] ^ d[38] ^ d[13] ^ d[31] ;
o[1] = d[23] ^ c[19] ^ c[12] ^ d[47] ^ d[40] ^ c[28] ^ c[21] ^ d[41] ^ c[0] ^ c[30] ^ d[10] ^ c[22] ^ c[8] ^ c[1] ^ d[34] ^ d[0] ^ c[31] ^ d[35] ^ d[1] ^ d[20] ^ d[19] ^ d[12] ^ d[9] ^ d[36] ^ d[13] ^ c[17] ^ d[3] ^ d[30] ^ d[14] ^ c[18] ^ c[11] ^ d[46] ^ d[38] ^ d[31] ;
o[2] = d[23] ^ d[15] ^ c[20] ^ c[19] ^ d[47] ^ d[40] ^ d[39] ^ c[28] ^ d[16] ^ c[21] ^ d[41] ^ c[0] ^ d[33] ^ d[17] ^ d[10] ^ c[22] ^ c[14] ^ c[8] ^ c[1] ^ d[34] ^ d[11] ^ c[23] ^ c[15] ^ c[2] ^ d[8] ^ d[12] ^ c[16] ^ d[9] ^ d[21] ^ c[10] ^ d[45] ^ d[29] ^ d[3] ^ d[30] ^ d[46] ^ d[38] ^ d[31] ;
o[3] = d[15] ^ c[20] ^ d[40] ^ d[39] ^ d[32] ^ d[16] ^ c[21] ^ d[33] ^ c[29] ^ d[10] ^ c[22] ^ c[1] ^ d[7] ^ c[23] ^ d[11] ^ c[15] ^ c[9] ^ c[2] ^ d[8] ^ d[20] ^ c[24] ^ c[16] ^ c[3] ^ d[44] ^ d[9] ^ d[28] ^ d[2] ^ c[17] ^ d[45] ^ d[37] ^ d[30] ^ d[29] ^ d[22] ^ d[14] ^ c[11] ^ d[46] ^ d[38] ;
o[4] = d[23] ^ d[47] ^ d[39] ^ d[32] ^ c[28] ^ d[16] ^ c[13] ^ d[41] ^ d[6] ^ d[17] ^ c[29] ^ c[30] ^ c[22] ^ c[14] ^ c[8] ^ d[7] ^ d[0] ^ c[31] ^ d[18] ^ c[23] ^ c[15] ^ c[9] ^ c[2] ^ d[43] ^ d[35] ^ d[8] ^ d[1] ^ d[27] ^ c[24] ^ c[3] ^ d[44] ^ d[9] ^ d[36] ^ d[2] ^ d[28] ^ c[25] ^ c[17] ^ c[4] ^ d[45] ^ d[29] ^ d[3] ^ d[22] ^ d[14] ;
o[5] = d[23] ^ c[12] ^ d[47] ^ d[40] ^ d[5] ^ c[28] ^ c[21] ^ c[13] ^ d[41] ^ d[6] ^ c[30] ^ d[10] ^ c[8] ^ d[42] ^ d[7] ^ d[34] ^ d[26] ^ d[18] ^ c[23] ^ d[43] ^ d[8] ^ d[1] ^ d[27] ^ d[19] ^ c[24] ^ c[3] ^ d[44] ^ d[28] ^ c[25] ^ c[4] ^ d[37] ^ d[3] ^ c[26] ^ c[5] ^ d[46] ;
o[6] = c[27] ^ c[6] ^ d[40] ^ d[39] ^ d[5] ^ c[13] ^ d[41] ^ d[6] ^ d[33] ^ d[25] ^ c[29] ^ d[17] ^ c[22] ^ c[14] ^ d[42] ^ d[7] ^ d[0] ^ d[26] ^ c[31] ^ d[18] ^ c[9] ^ d[43] ^ d[27] ^ c[24] ^ d[9] ^ d[36] ^ d[2] ^ c[25] ^ c[4] ^ d[45] ^ d[22] ^ c[26] ^ d[46] ^ c[5] ^ d[4] ;
o[7] = d[23] ^ c[27] ^ d[15] ^ c[12] ^ d[47] ^ c[6] ^ d[39] ^ d[40] ^ d[5] ^ d[32] ^ d[24] ^ c[21] ^ c[13] ^ c[7] ^ c[0] ^ d[6] ^ d[25] ^ c[29] ^ c[30] ^ d[10] ^ c[8] ^ d[42] ^ d[0] ^ d[26] ^ c[31] ^ d[18] ^ c[23] ^ c[9] ^ d[8] ^ d[1] ^ d[19] ^ c[16] ^ d[44] ^ d[2] ^ d[13] ^ c[25] ^ d[45] ^ d[37] ^ d[22] ^ c[26] ^ c[18] ^ c[5] ^ d[4] ^ d[31] ;
o[8] = c[27] ^ d[15] ^ c[19] ^ c[12] ^ d[47] ^ c[6] ^ d[39] ^ d[5] ^ d[24] ^ d[16] ^ c[21] ^ c[7] ^ d[25] ^ c[29] ^ c[30] ^ d[10] ^ c[22] ^ c[1] ^ d[7] ^ c[15] ^ d[43] ^ d[35] ^ d[1] ^ d[19] ^ c[24] ^ d[12] ^ c[16] ^ d[44] ^ d[9] ^ d[36] ^ d[2] ^ d[13] ^ c[17] ^ d[37] ^ d[30] ^ c[26] ^ d[14] ^ c[18] ^ d[46] ^ d[4] ;
o[9] = d[23] ^ c[27] ^ d[15] ^ c[19] ^ c[20] ^ d[24] ^ c[28] ^ c[13] ^ c[7] ^ d[6] ^ c[30] ^ c[22] ^ c[8] ^ d[42] ^ d[34] ^ d[0] ^ c[31] ^ d[18] ^ c[23] ^ d[11] ^ c[2] ^ d[43] ^ d[8] ^ d[35] ^ d[1] ^ d[12] ^ c[16] ^ d[9] ^ d[36] ^ c[25] ^ d[13] ^ c[17] ^ d[45] ^ d[3] ^ d[29] ^ d[14] ^ c[18] ^ d[46] ^ d[38] ^ d[4] ;
o[10] = d[15] ^ c[20] ^ c[19] ^ c[12] ^ d[47] ^ d[5] ^ d[16] ^ c[13] ^ c[0] ^ d[33] ^ d[42] ^ d[7] ^ d[34] ^ d[18] ^ d[11] ^ c[23] ^ c[15] ^ d[8] ^ d[19] ^ c[24] ^ d[12] ^ c[16] ^ c[3] ^ d[44] ^ d[28] ^ d[21] ^ c[17] ^ c[10] ^ d[45] ^ c[26] ^ d[14] ^ d[38] ^ d[31] ;
o[11] = d[23] ^ c[27] ^ c[20] ^ c[12] ^ d[47] ^ d[32] ^ c[28] ^ d[16] ^ c[0] ^ d[6] ^ d[33] ^ c[29] ^ c[8] ^ c[1] ^ d[7] ^ d[0] ^ c[31] ^ d[11] ^ c[15] ^ c[9] ^ d[43] ^ d[35] ^ d[27] ^ d[20] ^ d[19] ^ c[24] ^ d[44] ^ d[2] ^ d[21] ^ c[25] ^ c[17] ^ c[10] ^ c[4] ^ d[3] ^ d[30] ^ d[22] ^ d[14] ^ c[11] ^ d[46] ^ d[38] ^ d[4] ^ d[31] ;
o[12] = d[23] ^ d[47] ^ d[5] ^ d[32] ^ d[16] ^ d[41] ^ d[6] ^ d[17] ^ c[30] ^ c[14] ^ c[8] ^ c[1] ^ d[42] ^ d[34] ^ d[0] ^ d[26] ^ c[31] ^ c[15] ^ c[2] ^ d[43] ^ d[35] ^ d[1] ^ d[20] ^ c[25] ^ d[45] ^ d[29] ^ d[30] ^ c[26] ^ c[11] ^ c[5] ^ d[46] ^ d[38] ;
o[13] = c[27] ^ d[15] ^ c[12] ^ c[6] ^ d[40] ^ d[5] ^ d[16] ^ c[0] ^ d[41] ^ d[33] ^ d[25] ^ d[42] ^ d[34] ^ d[0] ^ c[31] ^ c[15] ^ c[9] ^ c[2] ^ d[19] ^ c[16] ^ c[3] ^ d[44] ^ d[28] ^ d[45] ^ d[37] ^ d[29] ^ d[22] ^ c[26] ^ d[46] ^ d[4] ^ d[31] ;
o[14] = d[15] ^ c[27] ^ d[39] ^ d[40] ^ d[32] ^ d[24] ^ c[28] ^ c[13] ^ c[7] ^ d[41] ^ d[33] ^ c[1] ^ d[18] ^ d[43] ^ d[27] ^ c[16] ^ d[44] ^ c[3] ^ d[36] ^ d[28] ^ d[21] ^ c[17] ^ c[10] ^ d[45] ^ c[4] ^ d[3] ^ d[30] ^ d[14] ^ d[4] ;
o[15] = d[23] ^ d[40] ^ d[39] ^ d[32] ^ c[28] ^ c[0] ^ c[29] ^ d[17] ^ c[14] ^ c[8] ^ d[42] ^ d[26] ^ c[2] ^ d[43] ^ d[35] ^ d[27] ^ d[20] ^ d[44] ^ d[2] ^ d[13] ^ c[17] ^ c[4] ^ d[3] ^ d[29] ^ d[14] ^ c[18] ^ c[11] ^ c[5] ^ d[38] ^ d[31] ;
o[16] = d[23] ^ d[15] ^ c[19] ^ d[47] ^ c[6] ^ d[39] ^ c[28] ^ c[21] ^ c[13] ^ d[25] ^ d[17] ^ c[30] ^ d[10] ^ c[14] ^ c[8] ^ d[42] ^ c[1] ^ d[34] ^ d[0] ^ d[26] ^ c[31] ^ d[18] ^ d[43] ^ d[35] ^ d[1] ^ d[12] ^ c[16] ^ c[3] ^ d[28] ^ d[21] ^ c[10] ^ d[3] ^ d[30] ^ c[5] ;
o[17] = c[20] ^ c[6] ^ d[24] ^ d[16] ^ c[7] ^ d[41] ^ d[33] ^ d[25] ^ c[29] ^ d[17] ^ c[22] ^ c[14] ^ d[42] ^ d[34] ^ d[0] ^ c[31] ^ d[11] ^ c[15] ^ c[9] ^ c[2] ^ d[27] ^ d[20] ^ d[9] ^ d[2] ^ c[17] ^ c[4] ^ d[29] ^ d[22] ^ d[14] ^ c[11] ^ d[46] ^ d[38] ;
o[18] = d[23] ^ d[15] ^ c[12] ^ d[40] ^ d[32] ^ d[24] ^ d[16] ^ c[21] ^ c[7] ^ d[41] ^ d[33] ^ c[30] ^ d[10] ^ c[8] ^ d[26] ^ c[23] ^ c[15] ^ d[8] ^ d[1] ^ d[19] ^ c[16] ^ c[3] ^ d[28] ^ d[21] ^ d[13] ^ c[10] ^ d[45] ^ d[37] ^ c[18] ^ c[5] ;
o[19] = d[23] ^ d[15] ^ c[19] ^ c[6] ^ d[39] ^ d[40] ^ d[32] ^ c[13] ^ c[0] ^ d[25] ^ c[22] ^ c[8] ^ d[7] ^ d[0] ^ c[31] ^ d[18] ^ c[9] ^ d[27] ^ d[20] ^ c[24] ^ d[12] ^ c[16] ^ d[44] ^ d[9] ^ d[36] ^ c[17] ^ c[4] ^ d[22] ^ d[14] ^ c[11] ^ d[31] ;
o[20] = c[20] ^ c[12] ^ d[39] ^ d[24] ^ c[7] ^ c[0] ^ d[6] ^ d[17] ^ c[14] ^ c[1] ^ d[26] ^ d[11] ^ c[23] ^ c[9] ^ d[43] ^ d[8] ^ d[35] ^ d[19] ^ d[21] ^ d[13] ^ c[25] ^ c[17] ^ c[10] ^ d[30] ^ d[22] ^ d[14] ^ c[18] ^ c[5] ^ d[38] ^ d[31] ;
o[21] = d[23] ^ c[19] ^ c[6] ^ d[5] ^ d[16] ^ c[21] ^ c[13] ^ d[25] ^ d[10] ^ c[8] ^ d[42] ^ c[1] ^ d[7] ^ d[34] ^ d[18] ^ c[15] ^ c[2] ^ d[20] ^ d[12] ^ c[24] ^ d[21] ^ d[13] ^ c[10] ^ d[37] ^ d[30] ^ d[29] ^ c[26] ^ c[18] ^ c[11] ^ d[38] ;
o[22] = d[23] ^ c[27] ^ c[20] ^ c[19] ^ d[47] ^ d[24] ^ c[28] ^ d[16] ^ c[21] ^ c[13] ^ c[7] ^ c[0] ^ d[6] ^ d[33] ^ c[29] ^ d[10] ^ c[22] ^ c[8] ^ d[0] ^ c[31] ^ d[18] ^ d[11] ^ c[15] ^ c[2] ^ d[35] ^ d[20] ^ d[12] ^ c[3] ^ d[9] ^ d[36] ^ d[2] ^ d[28] ^ d[21] ^ d[13] ^ c[25] ^ c[10] ^ d[29] ^ d[3] ^ c[18] ^ c[11] ^ d[38] ^ d[4] ^ d[31] ;
o[23] = c[20] ^ c[19] ^ d[47] ^ d[5] ^ d[32] ^ d[16] ^ c[13] ^ d[41] ^ c[0] ^ c[30] ^ c[22] ^ c[1] ^ d[34] ^ d[0] ^ c[31] ^ d[18] ^ d[11] ^ c[23] ^ c[15] ^ d[8] ^ d[1] ^ d[27] ^ d[20] ^ d[12] ^ c[3] ^ d[9] ^ d[28] ^ d[21] ^ d[13] ^ c[10] ^ c[4] ^ d[30] ^ c[26] ^ c[18] ^ c[11] ^ d[46] ^ d[38] ^ d[31] ;
o[24] = c[27] ^ d[15] ^ c[19] ^ c[20] ^ c[12] ^ d[40] ^ c[21] ^ c[0] ^ d[33] ^ d[17] ^ d[10] ^ c[14] ^ c[1] ^ d[7] ^ d[0] ^ d[26] ^ c[31] ^ c[23] ^ d[11] ^ c[2] ^ d[8] ^ d[27] ^ d[19] ^ d[20] ^ c[24] ^ d[12] ^ c[16] ^ c[4] ^ d[45] ^ d[37] ^ d[30] ^ d[29] ^ c[11] ^ d[46] ^ c[5] ^ d[4] ^ d[31] ;
o[25] = c[20] ^ c[12] ^ c[6] ^ d[39] ^ d[32] ^ c[28] ^ d[16] ^ c[21] ^ c[13] ^ d[6] ^ d[25] ^ c[22] ^ d[10] ^ c[1] ^ d[7] ^ d[26] ^ d[18] ^ d[11] ^ c[15] ^ c[2] ^ d[19] ^ c[24] ^ d[44] ^ c[3] ^ d[9] ^ d[36] ^ d[28] ^ c[25] ^ c[17] ^ d[45] ^ d[3] ^ d[30] ^ d[29] ^ d[14] ^ c[5] ;
o[26] = d[23] ^ c[12] ^ d[47] ^ c[6] ^ d[5] ^ d[24] ^ c[28] ^ d[16] ^ c[7] ^ d[41] ^ d[6] ^ d[25] ^ c[22] ^ c[8] ^ d[0] ^ c[31] ^ c[23] ^ c[15] ^ c[9] ^ c[2] ^ d[43] ^ d[8] ^ d[27] ^ d[19] ^ c[3] ^ d[44] ^ d[9] ^ d[28] ^ d[21] ^ c[25] ^ c[10] ^ c[4] ^ d[37] ^ d[29] ^ d[3] ^ d[22] ^ c[26] ;
o[27] = d[23] ^ c[27] ^ d[15] ^ d[40] ^ d[5] ^ d[24] ^ c[13] ^ c[7] ^ c[29] ^ c[8] ^ d[42] ^ d[7] ^ d[26] ^ d[18] ^ c[23] ^ c[9] ^ d[43] ^ d[8] ^ d[27] ^ d[20] ^ c[24] ^ c[16] ^ c[3] ^ d[36] ^ d[28] ^ d[2] ^ d[21] ^ c[10] ^ c[4] ^ d[22] ^ c[26] ^ c[11] ^ d[46] ^ c[5] ^ d[4] ;
o[28] = d[23] ^ c[27] ^ c[12] ^ c[6] ^ d[39] ^ c[28] ^ d[41] ^ d[6] ^ d[25] ^ c[30] ^ d[17] ^ c[14] ^ c[8] ^ d[42] ^ d[7] ^ d[26] ^ c[9] ^ d[35] ^ d[27] ^ d[1] ^ d[20] ^ d[19] ^ c[24] ^ d[21] ^ c[25] ^ c[17] ^ c[10] ^ d[45] ^ c[4] ^ d[3] ^ d[22] ^ d[14] ^ c[11] ^ c[5] ^ d[4] ;
o[29] = c[12] ^ c[6] ^ d[40] ^ d[5] ^ d[24] ^ d[16] ^ c[28] ^ c[13] ^ c[7] ^ d[41] ^ d[6] ^ d[25] ^ c[29] ^ d[34] ^ d[26] ^ d[0] ^ c[31] ^ d[18] ^ c[15] ^ c[9] ^ d[20] ^ d[19] ^ d[44] ^ d[2] ^ d[21] ^ c[25] ^ d[13] ^ c[10] ^ d[3] ^ d[22] ^ c[26] ^ c[18] ^ c[11] ^ c[5] ^ d[38] ;
o[30] = d[23] ^ c[27] ^ d[15] ^ c[19] ^ c[12] ^ c[6] ^ d[40] ^ d[39] ^ d[5] ^ d[24] ^ c[13] ^ c[7] ^ d[33] ^ d[25] ^ c[30] ^ c[29] ^ d[17] ^ c[14] ^ c[8] ^ d[18] ^ d[43] ^ d[1] ^ d[19] ^ d[20] ^ d[12] ^ c[16] ^ d[2] ^ d[21] ^ c[10] ^ d[37] ^ c[26] ^ c[11] ^ d[4] ;
o[31] = c[17] ^ d[23] ^ c[27] ^ c[9] ^ c[20] ^ c[30] ^ d[17] ^ c[12] ^ d[1] ^ d[20] ^ c[14] ^ d[19] ^ d[3] ^ d[22] ^ d[39] ^ d[14] ^ c[8] ^ d[32] ^ d[42] ^ d[24] ^ c[28] ^ c[11] ^ d[16] ^ d[0] ^ d[36] ^ d[18] ^ c[31] ^ c[13] ^ d[11] ^ c[15] ^ d[38] ^ d[4] ^ c[7] ;
        crc6B = o;
    end
    endfunction // crc6B

    ////////////////////////////////////////////////
    // crc5B
    ////////////////////////////////////////////////
    function [31:0] crc5B (
        input        [31:0]      c,
        input        [39:0]      d
        );
    reg          [31:0]      o;
    begin
o[0] = c[17] ^ d[23] ^ d[33] ^ d[15] ^ c[20] ^ c[2] ^ c[29] ^ d[8] ^ d[27] ^ c[22] ^ c[4] ^ d[10] ^ c[24] ^ d[30] ^ d[29] ^ d[39] ^ c[16] ^ d[5] ^ c[26] ^ d[14] ^ c[8] ^ c[18] ^ c[1] ^ d[7] ^ c[21] ^ d[9] ^ d[2] ^ d[11] ^ c[23] ^ d[13] ;
o[1] = d[23] ^ d[33] ^ d[15] ^ d[6] ^ c[27] ^ c[9] ^ c[19] ^ c[20] ^ c[29] ^ c[30] ^ d[27] ^ d[1] ^ c[4] ^ d[12] ^ d[30] ^ d[39] ^ c[16] ^ d[22] ^ d[5] ^ c[26] ^ c[8] ^ d[32] ^ c[1] ^ d[26] ^ c[3] ^ d[2] ^ d[11] ^ c[5] ^ d[28] ^ d[38] ^ c[25] ^ d[4] ;
o[2] = d[23] ^ c[0] ^ d[33] ^ d[15] ^ c[10] ^ c[27] ^ c[9] ^ d[25] ^ c[29] ^ c[30] ^ d[8] ^ c[22] ^ d[1] ^ d[37] ^ d[3] ^ c[24] ^ d[30] ^ c[6] ^ d[39] ^ c[16] ^ d[22] ^ c[8] ^ d[32] ^ c[18] ^ c[1] ^ c[28] ^ d[7] ^ d[0] ^ d[26] ^ d[9] ^ c[31] ^ d[2] ^ c[23] ^ c[5] ^ d[21] ^ d[38] ^ d[4] ^ d[13] ^ d[31] ;
o[3] = c[17] ^ c[0] ^ d[6] ^ c[9] ^ c[10] ^ c[19] ^ c[2] ^ d[25] ^ d[8] ^ c[29] ^ c[30] ^ d[1] ^ d[20] ^ d[37] ^ c[24] ^ d[3] ^ d[12] ^ d[29] ^ c[6] ^ d[30] ^ d[22] ^ d[32] ^ d[14] ^ d[24] ^ c[1] ^ c[11] ^ d[7] ^ c[28] ^ d[0] ^ c[31] ^ d[36] ^ d[2] ^ c[23] ^ d[38] ^ d[21] ^ c[25] ^ d[31] ^ c[7] ;
o[4] = d[15] ^ c[12] ^ d[39] ^ d[24] ^ c[21] ^ c[7] ^ c[0] ^ d[33] ^ d[6] ^ c[30] ^ c[22] ^ d[10] ^ d[0] ^ c[31] ^ c[23] ^ d[8] ^ d[35] ^ d[27] ^ d[1] ^ d[20] ^ d[19] ^ c[16] ^ c[3] ^ d[9] ^ d[36] ^ d[28] ^ d[21] ^ c[25] ^ c[17] ^ c[10] ^ c[4] ^ d[37] ^ d[14] ^ c[11] ^ d[31] ;
o[5] = d[15] ^ c[20] ^ c[12] ^ d[39] ^ d[32] ^ c[21] ^ c[13] ^ d[33] ^ c[29] ^ d[10] ^ d[34] ^ d[0] ^ d[26] ^ c[31] ^ d[18] ^ d[11] ^ c[2] ^ d[35] ^ d[20] ^ d[19] ^ c[16] ^ d[36] ^ d[2] ^ d[29] ^ c[11] ^ c[5] ^ d[38] ;
o[6] = c[12] ^ c[6] ^ d[32] ^ c[21] ^ c[13] ^ c[0] ^ d[33] ^ d[25] ^ c[30] ^ d[17] ^ d[10] ^ c[22] ^ c[14] ^ d[34] ^ d[18] ^ d[35] ^ d[1] ^ d[19] ^ c[3] ^ d[9] ^ d[28] ^ c[17] ^ d[37] ^ d[14] ^ d[38] ^ d[31] ;
o[7] = d[23] ^ d[15] ^ c[20] ^ d[39] ^ d[5] ^ d[32] ^ d[24] ^ d[16] ^ c[21] ^ c[13] ^ c[7] ^ c[0] ^ c[29] ^ d[17] ^ d[10] ^ c[14] ^ c[8] ^ d[7] ^ d[34] ^ d[0] ^ c[31] ^ d[18] ^ d[11] ^ c[15] ^ c[2] ^ c[24] ^ c[16] ^ d[36] ^ d[2] ^ c[17] ^ d[37] ^ d[29] ^ c[26] ^ d[14] ^ d[31] ;
o[8] = c[0] ^ d[6] ^ c[27] ^ c[9] ^ c[20] ^ c[2] ^ c[29] ^ c[30] ^ d[8] ^ d[17] ^ d[35] ^ d[27] ^ d[1] ^ c[4] ^ c[14] ^ c[24] ^ d[29] ^ d[39] ^ d[22] ^ d[5] ^ c[26] ^ d[7] ^ d[16] ^ c[3] ^ d[36] ^ d[2] ^ d[11] ^ c[23] ^ d[28] ^ d[38] ^ c[15] ^ c[25] ^ d[4] ^ d[31] ;
o[9] = c[27] ^ d[6] ^ d[15] ^ c[10] ^ c[30] ^ d[35] ^ d[1] ^ d[10] ^ d[27] ^ c[4] ^ d[37] ^ c[24] ^ d[3] ^ d[30] ^ c[16] ^ d[5] ^ c[26] ^ c[1] ^ d[7] ^ d[16] ^ c[28] ^ d[34] ^ d[26] ^ d[0] ^ c[21] ^ c[3] ^ c[31] ^ c[5] ^ d[28] ^ d[38] ^ c[15] ^ d[21] ^ d[4] ^ c[25] ;
o[10] = d[23] ^ c[27] ^ c[20] ^ c[6] ^ d[39] ^ c[28] ^ c[21] ^ d[6] ^ d[25] ^ d[10] ^ c[8] ^ c[1] ^ d[7] ^ d[34] ^ d[0] ^ d[26] ^ c[31] ^ d[11] ^ c[23] ^ d[8] ^ d[20] ^ c[24] ^ d[36] ^ c[25] ^ d[13] ^ d[37] ^ d[3] ^ d[30] ^ c[18] ^ c[11] ^ c[5] ^ d[4] ;
o[11] = c[17] ^ d[23] ^ d[15] ^ d[6] ^ c[9] ^ c[19] ^ c[20] ^ d[25] ^ d[8] ^ c[12] ^ d[35] ^ d[27] ^ c[4] ^ d[19] ^ d[3] ^ d[12] ^ d[30] ^ c[6] ^ d[39] ^ c[16] ^ d[22] ^ d[14] ^ c[8] ^ d[24] ^ c[18] ^ c[1] ^ c[28] ^ d[36] ^ d[11] ^ c[23] ^ d[38] ^ c[25] ^ c[7] ^ d[13] ;
o[12] = d[33] ^ d[15] ^ c[10] ^ c[9] ^ c[19] ^ d[8] ^ d[35] ^ d[27] ^ c[22] ^ c[4] ^ d[37] ^ d[12] ^ d[30] ^ d[39] ^ c[16] ^ d[22] ^ d[24] ^ c[1] ^ d[34] ^ d[26] ^ d[9] ^ d[18] ^ c[13] ^ c[23] ^ c[5] ^ d[21] ^ d[38] ^ c[7] ;
o[13] = c[17] ^ d[23] ^ c[10] ^ d[33] ^ c[20] ^ c[2] ^ d[25] ^ d[8] ^ d[17] ^ d[20] ^ c[14] ^ d[37] ^ c[24] ^ d[29] ^ c[6] ^ d[32] ^ d[14] ^ c[8] ^ c[11] ^ d[7] ^ d[34] ^ d[26] ^ d[36] ^ c[23] ^ d[11] ^ c[5] ^ d[38] ^ d[21] ;
o[14] = c[0] ^ d[6] ^ c[9] ^ d[33] ^ d[25] ^ c[12] ^ d[35] ^ d[10] ^ d[37] ^ d[19] ^ d[20] ^ c[24] ^ c[6] ^ d[22] ^ d[32] ^ c[18] ^ d[24] ^ d[7] ^ d[16] ^ c[11] ^ c[21] ^ c[3] ^ d[36] ^ d[28] ^ c[15] ^ d[31] ^ d[13] ^ c[25] ^ c[7] ;
o[15] = d[23] ^ c[0] ^ d[6] ^ d[15] ^ c[10] ^ c[19] ^ d[35] ^ c[12] ^ c[22] ^ d[27] ^ c[4] ^ d[19] ^ d[30] ^ d[12] ^ c[16] ^ d[5] ^ c[26] ^ c[8] ^ d[32] ^ d[24] ^ c[1] ^ d[34] ^ d[36] ^ d[18] ^ d[9] ^ c[13] ^ d[21] ^ c[25] ^ c[7] ^ d[31] ;
o[16] = d[15] ^ c[27] ^ d[39] ^ c[21] ^ c[13] ^ c[0] ^ c[29] ^ d[17] ^ c[22] ^ d[10] ^ c[14] ^ d[7] ^ d[34] ^ d[26] ^ d[18] ^ c[9] ^ d[35] ^ d[27] ^ d[20] ^ c[24] ^ c[16] ^ d[9] ^ d[2] ^ d[13] ^ c[4] ^ d[22] ^ c[18] ^ c[11] ^ c[5] ^ d[4] ^ d[31] ;
o[17] = c[17] ^ d[6] ^ d[33] ^ c[10] ^ c[19] ^ d[25] ^ d[8] ^ c[30] ^ d[17] ^ c[12] ^ d[1] ^ c[22] ^ c[14] ^ d[19] ^ d[3] ^ d[12] ^ c[6] ^ d[30] ^ d[14] ^ c[1] ^ d[16] ^ c[28] ^ d[34] ^ d[26] ^ d[9] ^ c[23] ^ c[5] ^ d[38] ^ c[15] ^ d[21] ^ c[25] ;
o[18] = d[15] ^ d[33] ^ d[25] ^ c[20] ^ c[2] ^ c[29] ^ d[8] ^ d[37] ^ d[20] ^ c[24] ^ c[6] ^ d[29] ^ c[16] ^ d[5] ^ c[26] ^ d[32] ^ c[18] ^ d[24] ^ d[7] ^ d[16] ^ c[11] ^ d[0] ^ c[31] ^ d[18] ^ c[13] ^ d[2] ^ d[11] ^ c[23] ^ c[15] ^ d[13] ^ c[7] ;
o[19] = c[17] ^ d[23] ^ c[0] ^ d[6] ^ d[15] ^ c[27] ^ c[19] ^ c[30] ^ d[17] ^ c[12] ^ d[1] ^ d[10] ^ c[14] ^ d[19] ^ d[12] ^ c[24] ^ c[16] ^ d[14] ^ d[32] ^ c[8] ^ d[24] ^ d[7] ^ c[21] ^ c[3] ^ d[36] ^ d[28] ^ c[25] ^ d[4] ^ c[7] ^ d[31] ;
o[20] = d[23] ^ c[17] ^ c[0] ^ d[6] ^ c[9] ^ c[20] ^ d[35] ^ c[22] ^ d[27] ^ c[4] ^ d[3] ^ d[30] ^ d[22] ^ d[5] ^ c[26] ^ d[14] ^ c[8] ^ c[18] ^ c[1] ^ c[28] ^ d[16] ^ d[0] ^ c[31] ^ d[9] ^ d[18] ^ c[13] ^ d[11] ^ c[15] ^ d[13] ^ c[25] ^ d[31] ;
o[21] = c[27] ^ c[9] ^ d[15] ^ c[10] ^ c[19] ^ c[2] ^ c[29] ^ d[8] ^ d[17] ^ d[10] ^ c[14] ^ d[12] ^ d[30] ^ d[29] ^ d[22] ^ c[16] ^ d[5] ^ c[26] ^ c[18] ^ c[1] ^ d[34] ^ c[21] ^ d[26] ^ d[2] ^ c[23] ^ c[5] ^ d[21] ^ d[4] ^ d[13] ;
o[22] = d[23] ^ d[15] ^ c[10] ^ c[27] ^ c[19] ^ d[25] ^ c[29] ^ c[30] ^ d[8] ^ d[27] ^ d[1] ^ c[4] ^ d[10] ^ d[20] ^ d[3] ^ d[12] ^ d[30] ^ c[6] ^ d[39] ^ c[16] ^ d[5] ^ c[26] ^ c[8] ^ c[18] ^ c[1] ^ c[28] ^ c[11] ^ d[16] ^ c[21] ^ c[3] ^ d[2] ^ c[23] ^ d[28] ^ d[21] ^ c[15] ^ d[4] ^ d[13] ;
o[23] = d[23] ^ d[33] ^ c[27] ^ c[9] ^ c[19] ^ c[30] ^ d[8] ^ c[12] ^ d[1] ^ d[10] ^ d[20] ^ d[19] ^ d[3] ^ d[12] ^ d[30] ^ d[39] ^ d[22] ^ d[5] ^ c[26] ^ c[8] ^ d[24] ^ c[18] ^ c[1] ^ c[28] ^ c[11] ^ d[0] ^ c[21] ^ d[26] ^ c[31] ^ c[23] ^ c[5] ^ d[38] ^ d[4] ^ c[7] ^ d[13] ;
o[24] = d[23] ^ c[27] ^ c[9] ^ c[10] ^ c[20] ^ c[19] ^ c[2] ^ d[25] ^ c[29] ^ c[12] ^ c[22] ^ d[19] ^ d[37] ^ c[24] ^ d[3] ^ d[12] ^ d[29] ^ c[6] ^ d[22] ^ d[32] ^ c[8] ^ d[7] ^ c[28] ^ d[0] ^ c[31] ^ d[9] ^ d[18] ^ c[13] ^ d[2] ^ d[11] ^ d[38] ^ d[21] ^ d[4] ;
o[25] = c[0] ^ d[6] ^ c[9] ^ c[10] ^ c[20] ^ c[30] ^ c[29] ^ d[8] ^ d[17] ^ d[1] ^ d[10] ^ d[37] ^ c[14] ^ d[20] ^ d[3] ^ d[22] ^ d[24] ^ c[28] ^ c[11] ^ c[21] ^ c[3] ^ d[18] ^ c[13] ^ d[36] ^ d[2] ^ d[11] ^ d[28] ^ c[23] ^ d[21] ^ d[31] ^ c[25] ^ c[7] ;
o[26] = c[17] ^ d[33] ^ d[15] ^ c[10] ^ c[20] ^ c[2] ^ c[30] ^ d[8] ^ d[17] ^ c[12] ^ d[35] ^ d[1] ^ c[14] ^ d[20] ^ d[19] ^ d[29] ^ d[39] ^ c[16] ^ d[14] ^ c[18] ^ c[11] ^ d[16] ^ d[0] ^ c[31] ^ d[36] ^ d[11] ^ c[23] ^ d[21] ^ c[15] ^ d[13] ;
o[27] = c[17] ^ d[15] ^ c[19] ^ c[12] ^ d[35] ^ d[10] ^ d[20] ^ d[19] ^ c[24] ^ d[12] ^ c[16] ^ d[32] ^ d[14] ^ c[18] ^ c[11] ^ d[7] ^ d[16] ^ d[34] ^ d[0] ^ c[21] ^ c[3] ^ c[31] ^ d[18] ^ c[13] ^ d[28] ^ d[38] ^ c[15] ^ d[13] ;
o[28] = c[0] ^ c[17] ^ d[6] ^ d[15] ^ d[33] ^ c[19] ^ c[20] ^ c[12] ^ d[17] ^ c[22] ^ d[27] ^ c[4] ^ d[37] ^ d[19] ^ c[14] ^ d[12] ^ c[16] ^ d[14] ^ c[18] ^ d[34] ^ d[9] ^ d[18] ^ c[13] ^ d[11] ^ d[31] ^ d[13] ^ c[25] ;
o[29] = c[17] ^ d[33] ^ c[19] ^ c[20] ^ d[8] ^ d[17] ^ d[10] ^ c[14] ^ d[30] ^ d[12] ^ d[5] ^ c[26] ^ d[14] ^ d[32] ^ c[1] ^ c[18] ^ d[16] ^ c[21] ^ d[26] ^ d[36] ^ d[18] ^ c[13] ^ c[23] ^ d[11] ^ c[5] ^ c[15] ^ d[13] ;
o[30] = c[0] ^ c[27] ^ d[15] ^ c[20] ^ c[2] ^ d[25] ^ c[19] ^ d[35] ^ d[17] ^ d[10] ^ c[22] ^ c[14] ^ d[29] ^ c[24] ^ c[6] ^ d[12] ^ c[16] ^ d[32] ^ c[18] ^ d[7] ^ d[16] ^ c[21] ^ d[9] ^ d[11] ^ c[15] ^ d[4] ^ d[13] ^ d[31] ;
o[31] = c[17] ^ c[0] ^ d[6] ^ d[15] ^ c[19] ^ c[20] ^ d[8] ^ d[10] ^ c[22] ^ d[3] ^ d[12] ^ d[30] ^ c[16] ^ d[14] ^ d[24] ^ c[1] ^ d[34] ^ d[16] ^ c[28] ^ c[21] ^ c[3] ^ d[9] ^ d[28] ^ c[23] ^ d[11] ^ c[15] ^ c[25] ^ c[7] ^ d[31] ;
        crc5B = o;
    end
    endfunction // crc5B

    ////////////////////////////////////////////////
    // crc4B
    ////////////////////////////////////////////////
    function [31:0] crc4B (
        input        [31:0]      c,
        input        [31:0]      d
        );
    reg          [31:0]      o;
    begin
o[0] = c[0] ^ d[6] ^ d[15] ^ c[9] ^ c[10] ^ d[25] ^ c[30] ^ c[12] ^ c[29] ^ d[1] ^ d[19] ^ c[24] ^ d[3] ^ c[6] ^ c[16] ^ d[22] ^ d[5] ^ c[26] ^ d[7] ^ c[28] ^ d[0] ^ c[31] ^ d[2] ^ d[21] ^ d[31] ^ c[25] ;
o[1] = c[0] ^ c[17] ^ c[27] ^ d[15] ^ c[9] ^ d[25] ^ c[12] ^ d[19] ^ d[20] ^ c[24] ^ d[3] ^ c[6] ^ d[30] ^ c[16] ^ d[22] ^ d[14] ^ d[24] ^ c[1] ^ d[7] ^ c[28] ^ c[11] ^ d[18] ^ c[13] ^ d[31] ^ d[4] ^ c[7] ;
o[2] = c[0] ^ c[17] ^ d[23] ^ d[15] ^ c[9] ^ d[25] ^ c[2] ^ c[30] ^ d[17] ^ d[1] ^ c[14] ^ c[24] ^ c[6] ^ d[30] ^ d[29] ^ c[16] ^ d[22] ^ d[5] ^ c[26] ^ d[14] ^ c[8] ^ c[18] ^ d[24] ^ c[1] ^ d[7] ^ d[0] ^ c[31] ^ d[18] ^ c[13] ^ d[31] ^ d[13] ^ c[7] ;
o[3] = c[17] ^ d[23] ^ d[6] ^ c[27] ^ c[10] ^ c[9] ^ c[19] ^ c[2] ^ d[17] ^ c[14] ^ d[30] ^ d[12] ^ d[29] ^ d[22] ^ d[14] ^ c[8] ^ d[24] ^ c[1] ^ c[18] ^ d[16] ^ d[0] ^ c[3] ^ c[31] ^ d[28] ^ d[21] ^ c[15] ^ c[25] ^ d[4] ^ c[7] ^ d[13] ;
o[4] = c[0] ^ d[23] ^ d[6] ^ d[25] ^ c[19] ^ c[20] ^ c[2] ^ c[30] ^ c[12] ^ c[29] ^ d[1] ^ d[27] ^ c[4] ^ d[19] ^ d[20] ^ c[24] ^ c[6] ^ d[12] ^ d[29] ^ c[8] ^ c[18] ^ d[7] ^ d[16] ^ c[11] ^ d[0] ^ c[3] ^ c[31] ^ d[2] ^ d[11] ^ d[28] ^ c[15] ^ d[31] ^ d[13] ^ c[25] ;
o[5] = c[0] ^ c[10] ^ d[25] ^ c[19] ^ c[20] ^ c[29] ^ d[10] ^ d[27] ^ c[4] ^ c[24] ^ d[3] ^ c[6] ^ d[12] ^ d[30] ^ d[24] ^ c[1] ^ d[7] ^ c[28] ^ c[21] ^ c[3] ^ d[26] ^ d[18] ^ c[13] ^ d[2] ^ d[11] ^ d[28] ^ c[5] ^ d[21] ^ d[31] ^ c[7] ;
o[6] = d[23] ^ d[6] ^ c[20] ^ c[2] ^ d[25] ^ c[29] ^ c[30] ^ d[17] ^ c[22] ^ d[1] ^ d[10] ^ d[27] ^ c[4] ^ d[20] ^ c[14] ^ d[30] ^ d[29] ^ c[6] ^ c[8] ^ d[24] ^ c[1] ^ c[11] ^ c[21] ^ d[26] ^ d[9] ^ d[2] ^ d[11] ^ c[5] ^ c[25] ^ c[7] ;
o[7] = c[0] ^ d[23] ^ d[6] ^ d[15] ^ c[10] ^ c[2] ^ c[29] ^ d[8] ^ d[10] ^ c[22] ^ c[24] ^ d[3] ^ d[29] ^ c[16] ^ c[8] ^ d[24] ^ d[7] ^ c[28] ^ d[16] ^ c[21] ^ c[3] ^ d[26] ^ d[9] ^ d[2] ^ c[23] ^ d[28] ^ c[5] ^ c[15] ^ d[21] ^ d[31] ^ c[25] ^ c[7] ;
o[8] = c[0] ^ c[17] ^ d[23] ^ c[10] ^ c[12] ^ d[8] ^ c[22] ^ d[27] ^ c[4] ^ d[19] ^ d[20] ^ d[3] ^ d[30] ^ d[14] ^ c[8] ^ c[1] ^ c[28] ^ c[11] ^ d[0] ^ c[3] ^ c[31] ^ d[9] ^ c[23] ^ d[28] ^ d[21] ^ d[31] ;
o[9] = c[9] ^ c[2] ^ c[29] ^ d[8] ^ c[12] ^ d[27] ^ c[4] ^ d[20] ^ d[19] ^ d[30] ^ d[29] ^ c[24] ^ d[22] ^ c[1] ^ c[18] ^ c[11] ^ d[7] ^ d[26] ^ d[18] ^ c[13] ^ d[2] ^ c[23] ^ c[5] ^ d[13] ;
o[10] = c[0] ^ d[15] ^ c[9] ^ c[19] ^ c[2] ^ c[29] ^ d[17] ^ c[14] ^ d[3] ^ d[12] ^ d[29] ^ c[16] ^ d[22] ^ d[5] ^ c[26] ^ c[28] ^ d[0] ^ c[3] ^ d[26] ^ c[31] ^ d[18] ^ c[13] ^ d[2] ^ d[28] ^ c[5] ^ d[31] ;
o[11] = c[0] ^ c[17] ^ c[27] ^ d[6] ^ d[15] ^ c[9] ^ c[20] ^ c[12] ^ d[17] ^ d[27] ^ c[4] ^ d[19] ^ c[14] ^ c[24] ^ d[3] ^ d[30] ^ c[16] ^ d[22] ^ d[5] ^ c[26] ^ d[14] ^ c[1] ^ d[7] ^ c[28] ^ d[16] ^ d[0] ^ c[3] ^ c[31] ^ d[11] ^ d[28] ^ c[15] ^ d[31] ^ d[4] ^ c[25] ;
o[12] = c[0] ^ c[17] ^ c[27] ^ c[9] ^ d[25] ^ c[2] ^ c[30] ^ c[12] ^ d[1] ^ d[10] ^ d[27] ^ c[4] ^ d[19] ^ c[24] ^ c[6] ^ d[30] ^ d[29] ^ d[22] ^ d[14] ^ c[18] ^ c[1] ^ d[7] ^ d[16] ^ d[0] ^ c[21] ^ d[26] ^ c[31] ^ d[18] ^ c[13] ^ c[5] ^ c[15] ^ d[31] ^ d[13] ^ d[4] ;
o[13] = d[6] ^ d[15] ^ c[10] ^ c[19] ^ c[2] ^ d[25] ^ d[17] ^ c[22] ^ c[14] ^ d[30] ^ d[12] ^ d[3] ^ d[29] ^ c[6] ^ c[16] ^ d[24] ^ c[1] ^ c[18] ^ c[28] ^ d[0] ^ c[3] ^ d[26] ^ d[18] ^ c[31] ^ d[9] ^ c[13] ^ d[28] ^ c[5] ^ d[21] ^ c[25] ^ c[7] ^ d[13] ;
o[14] = d[23] ^ c[17] ^ c[20] ^ c[2] ^ c[19] ^ d[25] ^ d[17] ^ c[29] ^ d[8] ^ d[27] ^ c[4] ^ c[14] ^ d[20] ^ d[29] ^ d[12] ^ c[6] ^ d[5] ^ c[26] ^ d[14] ^ c[8] ^ d[24] ^ c[11] ^ d[16] ^ c[3] ^ d[11] ^ d[2] ^ c[23] ^ d[28] ^ c[15] ^ c[7] ;
o[15] = d[23] ^ c[27] ^ c[9] ^ d[15] ^ c[20] ^ c[30] ^ c[12] ^ d[10] ^ d[1] ^ d[27] ^ c[4] ^ d[19] ^ c[24] ^ d[22] ^ c[16] ^ c[8] ^ c[18] ^ d[24] ^ d[16] ^ d[7] ^ c[21] ^ c[3] ^ d[26] ^ d[28] ^ d[11] ^ c[5] ^ c[15] ^ d[4] ^ d[13] ^ c[7] ;
o[16] = c[0] ^ c[17] ^ d[23] ^ c[19] ^ c[30] ^ c[12] ^ c[29] ^ d[1] ^ d[10] ^ c[22] ^ d[27] ^ c[4] ^ d[19] ^ c[24] ^ d[12] ^ d[5] ^ c[26] ^ d[14] ^ c[8] ^ d[7] ^ c[21] ^ d[26] ^ d[9] ^ d[18] ^ c[13] ^ d[2] ^ c[5] ^ d[31] ;
o[17] = d[6] ^ c[27] ^ c[9] ^ c[20] ^ d[25] ^ d[8] ^ c[30] ^ d[17] ^ c[22] ^ d[1] ^ c[14] ^ d[30] ^ c[6] ^ d[22] ^ c[1] ^ c[18] ^ d[0] ^ d[26] ^ d[18] ^ c[31] ^ d[9] ^ c[13] ^ c[23] ^ d[11] ^ c[5] ^ c[25] ^ d[4] ^ d[13] ;
o[18] = c[10] ^ c[2] ^ d[25] ^ c[19] ^ d[17] ^ d[8] ^ d[10] ^ c[14] ^ d[29] ^ c[24] ^ d[3] ^ c[6] ^ d[12] ^ d[5] ^ c[26] ^ d[24] ^ d[7] ^ c[28] ^ d[16] ^ d[0] ^ c[21] ^ c[31] ^ c[23] ^ c[15] ^ d[21] ^ c[7] ;
o[19] = d[23] ^ c[27] ^ d[6] ^ d[15] ^ c[20] ^ c[29] ^ c[22] ^ d[20] ^ c[24] ^ c[16] ^ c[8] ^ d[24] ^ d[16] ^ d[7] ^ c[11] ^ c[3] ^ d[9] ^ d[28] ^ d[2] ^ d[11] ^ c[15] ^ d[4] ^ c[25] ^ c[7] ;
o[20] = d[23] ^ c[17] ^ d[15] ^ d[6] ^ c[9] ^ c[30] ^ d[8] ^ c[12] ^ d[27] ^ d[1] ^ c[4] ^ d[10] ^ d[19] ^ d[3] ^ c[16] ^ d[22] ^ d[5] ^ c[26] ^ d[14] ^ c[8] ^ c[28] ^ c[21] ^ c[23] ^ c[25] ;
o[21] = c[17] ^ c[27] ^ c[9] ^ c[10] ^ c[29] ^ c[22] ^ c[24] ^ d[22] ^ d[14] ^ d[5] ^ c[26] ^ c[18] ^ d[7] ^ d[26] ^ d[0] ^ c[31] ^ d[9] ^ d[18] ^ c[13] ^ d[2] ^ c[5] ^ d[21] ^ d[4] ^ d[13] ;
o[22] = c[0] ^ c[27] ^ d[15] ^ c[9] ^ c[19] ^ c[12] ^ c[29] ^ d[8] ^ d[17] ^ d[19] ^ d[20] ^ c[14] ^ c[24] ^ d[12] ^ c[16] ^ d[22] ^ d[5] ^ c[26] ^ c[18] ^ d[7] ^ c[11] ^ d[0] ^ c[31] ^ d[2] ^ c[23] ^ d[31] ^ d[13] ^ d[4] ;
o[23] = c[0] ^ c[17] ^ c[27] ^ d[15] ^ c[9] ^ d[25] ^ c[19] ^ c[20] ^ c[29] ^ c[6] ^ d[12] ^ d[30] ^ c[16] ^ d[22] ^ d[5] ^ c[26] ^ d[14] ^ c[1] ^ d[16] ^ d[0] ^ c[31] ^ d[18] ^ c[13] ^ d[2] ^ d[11] ^ c[15] ^ d[31] ^ d[4] ;
o[24] = c[17] ^ d[15] ^ c[27] ^ c[10] ^ c[20] ^ c[2] ^ c[30] ^ d[17] ^ d[1] ^ d[10] ^ c[14] ^ d[30] ^ d[3] ^ d[29] ^ c[16] ^ d[14] ^ d[24] ^ c[1] ^ c[18] ^ c[28] ^ c[21] ^ d[11] ^ d[21] ^ d[4] ^ c[7] ^ d[13] ;
o[25] = d[23] ^ c[17] ^ c[2] ^ c[19] ^ c[29] ^ d[10] ^ c[22] ^ d[20] ^ d[29] ^ d[3] ^ d[12] ^ d[14] ^ c[8] ^ c[18] ^ c[28] ^ c[11] ^ d[16] ^ d[0] ^ c[21] ^ c[3] ^ c[31] ^ d[9] ^ d[2] ^ d[28] ^ c[15] ^ d[13] ;
o[26] = c[0] ^ d[6] ^ c[10] ^ d[25] ^ c[19] ^ c[20] ^ d[8] ^ c[22] ^ d[27] ^ c[4] ^ c[24] ^ d[3] ^ c[6] ^ d[12] ^ d[5] ^ c[26] ^ c[18] ^ d[7] ^ c[28] ^ d[0] ^ c[3] ^ c[31] ^ d[9] ^ d[11] ^ d[28] ^ c[23] ^ d[21] ^ d[31] ^ d[13] ^ c[25] ;
o[27] = d[6] ^ c[27] ^ c[19] ^ c[20] ^ c[29] ^ d[8] ^ d[10] ^ d[27] ^ c[4] ^ d[20] ^ d[30] ^ d[12] ^ c[24] ^ d[5] ^ c[26] ^ d[24] ^ c[1] ^ c[11] ^ d[7] ^ c[21] ^ d[26] ^ d[2] ^ c[23] ^ d[11] ^ c[5] ^ c[25] ^ d[4] ^ c[7] ;
o[28] = d[23] ^ c[27] ^ d[6] ^ c[20] ^ c[2] ^ d[25] ^ c[30] ^ c[12] ^ d[1] ^ d[10] ^ c[22] ^ d[19] ^ d[29] ^ c[24] ^ d[3] ^ c[6] ^ d[5] ^ c[26] ^ c[8] ^ d[7] ^ c[28] ^ c[21] ^ d[26] ^ d[9] ^ d[11] ^ c[5] ^ d[4] ^ c[25] ;
o[29] = c[27] ^ d[6] ^ c[9] ^ d[25] ^ c[29] ^ d[8] ^ d[10] ^ c[22] ^ d[3] ^ c[6] ^ d[22] ^ d[5] ^ c[26] ^ d[24] ^ c[28] ^ d[0] ^ c[21] ^ c[3] ^ c[31] ^ d[9] ^ d[18] ^ c[13] ^ d[28] ^ d[2] ^ c[23] ^ d[4] ^ c[25] ^ c[7] ;
o[30] = d[23] ^ c[10] ^ c[27] ^ c[29] ^ c[30] ^ d[8] ^ d[17] ^ d[27] ^ c[22] ^ d[1] ^ c[4] ^ c[14] ^ d[3] ^ c[24] ^ d[5] ^ c[26] ^ c[8] ^ d[24] ^ c[28] ^ d[7] ^ d[9] ^ d[2] ^ c[23] ^ d[21] ^ d[4] ^ c[7] ;
o[31] = d[23] ^ c[27] ^ d[6] ^ c[9] ^ d[8] ^ c[29] ^ c[30] ^ d[1] ^ d[20] ^ c[24] ^ d[3] ^ d[22] ^ c[8] ^ c[11] ^ d[7] ^ d[16] ^ c[28] ^ d[26] ^ d[0] ^ c[31] ^ d[2] ^ c[23] ^ c[5] ^ c[15] ^ d[4] ^ c[25] ;
        crc4B = o;
    end
    endfunction // crc4B

    ////////////////////////////////////////////////
    // crc3B
    ////////////////////////////////////////////////
    function [31:0] crc3B (
        input        [31:0]      c,
        input        [23:0]      d
        );
    reg          [31:0]      o;
    begin
o[0] = d[23] ^ c[17] ^ c[20] ^ d[17] ^ c[14] ^ c[24] ^ c[8] ^ d[14] ^ c[18] ^ d[7] ^ d[11] ^ d[13] ;
o[1] = d[23] ^ c[17] ^ d[6] ^ c[9] ^ c[20] ^ c[19] ^ d[17] ^ d[10] ^ c[14] ^ c[24] ^ d[12] ^ d[22] ^ d[14] ^ c[8] ^ d[7] ^ d[16] ^ c[21] ^ d[11] ^ c[15] ^ c[25] ;
o[2] = d[23] ^ c[17] ^ d[6] ^ c[9] ^ d[15] ^ c[10] ^ d[17] ^ d[10] ^ c[22] ^ c[14] ^ c[24] ^ d[22] ^ c[16] ^ d[5] ^ c[26] ^ d[14] ^ c[8] ^ d[7] ^ d[16] ^ c[21] ^ d[9] ^ c[15] ^ d[21] ^ c[25] ;
o[3] = c[17] ^ c[27] ^ d[6] ^ c[9] ^ d[15] ^ c[10] ^ d[8] ^ c[22] ^ d[20] ^ d[22] ^ c[16] ^ d[5] ^ c[26] ^ d[14] ^ c[18] ^ d[16] ^ c[11] ^ d[9] ^ c[23] ^ c[15] ^ d[21] ^ d[4] ^ c[25] ^ d[13] ;
o[4] = d[23] ^ c[27] ^ d[15] ^ c[10] ^ c[20] ^ c[19] ^ d[17] ^ d[8] ^ c[12] ^ c[14] ^ d[20] ^ d[19] ^ d[3] ^ d[12] ^ c[16] ^ d[5] ^ c[26] ^ c[8] ^ c[28] ^ c[11] ^ d[11] ^ c[23] ^ d[21] ^ d[4] ;
o[5] = d[23] ^ c[27] ^ c[9] ^ d[17] ^ c[29] ^ c[12] ^ d[10] ^ c[14] ^ d[20] ^ d[19] ^ d[3] ^ d[22] ^ c[8] ^ c[18] ^ c[28] ^ d[16] ^ c[11] ^ c[21] ^ d[18] ^ c[13] ^ d[2] ^ c[15] ^ d[4] ^ d[13] ;
o[6] = c[9] ^ d[15] ^ c[10] ^ c[19] ^ c[30] ^ c[29] ^ c[12] ^ d[17] ^ d[1] ^ c[22] ^ d[19] ^ c[14] ^ d[3] ^ d[12] ^ d[22] ^ c[16] ^ d[16] ^ c[28] ^ d[9] ^ d[18] ^ c[13] ^ d[2] ^ c[15] ^ d[21] ;
o[7] = d[23] ^ d[15] ^ c[10] ^ c[29] ^ c[30] ^ d[8] ^ d[1] ^ d[20] ^ c[24] ^ c[16] ^ c[8] ^ c[18] ^ d[7] ^ c[11] ^ d[16] ^ d[0] ^ c[31] ^ d[18] ^ c[13] ^ d[2] ^ c[23] ^ d[21] ^ c[15] ^ d[13] ;
o[8] = d[23] ^ d[6] ^ c[9] ^ d[15] ^ c[20] ^ c[19] ^ c[30] ^ c[12] ^ d[1] ^ d[20] ^ d[19] ^ d[12] ^ d[22] ^ c[16] ^ c[8] ^ c[18] ^ c[11] ^ d[0] ^ c[31] ^ d[11] ^ d[13] ^ c[25] ;
o[9] = c[17] ^ c[9] ^ c[10] ^ c[19] ^ c[20] ^ c[12] ^ d[10] ^ d[19] ^ d[12] ^ d[22] ^ d[5] ^ c[26] ^ d[14] ^ d[0] ^ c[21] ^ c[31] ^ d[18] ^ c[13] ^ d[11] ^ d[21] ;
o[10] = d[23] ^ c[17] ^ c[27] ^ c[10] ^ c[22] ^ d[10] ^ d[20] ^ c[24] ^ d[14] ^ c[8] ^ d[7] ^ c[11] ^ c[21] ^ d[9] ^ d[18] ^ c[13] ^ d[21] ^ d[4] ;
o[11] = d[23] ^ c[17] ^ d[6] ^ c[9] ^ c[20] ^ d[8] ^ c[12] ^ c[22] ^ d[20] ^ d[19] ^ c[24] ^ d[3] ^ d[22] ^ d[14] ^ c[8] ^ d[7] ^ c[28] ^ c[11] ^ d[9] ^ d[11] ^ c[23] ^ c[25] ;
o[12] = d[23] ^ c[17] ^ d[6] ^ c[9] ^ c[10] ^ c[20] ^ d[17] ^ c[29] ^ d[8] ^ c[12] ^ d[10] ^ c[14] ^ d[19] ^ d[22] ^ d[5] ^ c[26] ^ d[14] ^ c[8] ^ c[21] ^ d[18] ^ c[13] ^ d[11] ^ d[2] ^ c[23] ^ d[21] ^ c[25] ;
o[13] = c[27] ^ c[9] ^ c[10] ^ c[30] ^ d[17] ^ d[10] ^ d[1] ^ c[22] ^ d[20] ^ c[14] ^ c[24] ^ d[22] ^ d[5] ^ c[26] ^ c[18] ^ d[16] ^ d[7] ^ c[11] ^ c[21] ^ d[9] ^ d[18] ^ c[13] ^ c[15] ^ d[21] ^ d[4] ^ d[13] ;
o[14] = d[15] ^ d[6] ^ c[10] ^ c[27] ^ c[19] ^ d[8] ^ c[12] ^ d[17] ^ c[22] ^ d[20] ^ d[19] ^ c[14] ^ d[3] ^ d[12] ^ c[16] ^ c[28] ^ c[11] ^ d[16] ^ d[0] ^ d[9] ^ c[31] ^ c[23] ^ d[21] ^ c[15] ^ c[25] ^ d[4] ;
o[15] = c[17] ^ d[15] ^ c[20] ^ d[8] ^ c[29] ^ c[12] ^ d[20] ^ d[19] ^ c[24] ^ d[3] ^ c[16] ^ d[14] ^ d[5] ^ c[26] ^ c[11] ^ d[7] ^ c[28] ^ d[16] ^ d[18] ^ c[13] ^ d[2] ^ c[23] ^ d[11] ^ c[15] ;
o[16] = d[23] ^ c[27] ^ d[6] ^ d[15] ^ c[20] ^ c[29] ^ c[30] ^ c[12] ^ d[1] ^ d[10] ^ d[19] ^ c[16] ^ c[8] ^ c[21] ^ d[18] ^ c[13] ^ d[11] ^ d[2] ^ d[4] ^ c[25] ;
o[17] = c[17] ^ c[9] ^ c[30] ^ d[17] ^ d[10] ^ d[1] ^ c[22] ^ c[14] ^ d[3] ^ d[22] ^ d[5] ^ c[26] ^ d[14] ^ c[28] ^ d[0] ^ c[21] ^ c[31] ^ d[18] ^ d[9] ^ c[13] ;
o[18] = c[10] ^ c[27] ^ c[29] ^ d[17] ^ d[8] ^ c[22] ^ c[14] ^ c[18] ^ d[16] ^ d[0] ^ d[9] ^ c[31] ^ d[2] ^ c[23] ^ d[21] ^ c[15] ^ d[4] ^ d[13] ;
o[19] = d[15] ^ c[19] ^ d[8] ^ c[30] ^ d[1] ^ d[20] ^ c[24] ^ d[3] ^ d[12] ^ c[16] ^ c[11] ^ d[16] ^ d[7] ^ c[28] ^ c[23] ^ c[15] ;
o[20] = c[17] ^ d[15] ^ d[6] ^ c[20] ^ c[12] ^ c[29] ^ d[19] ^ c[24] ^ c[16] ^ d[14] ^ d[7] ^ d[0] ^ c[31] ^ d[2] ^ d[11] ^ c[25] ;
o[21] = c[17] ^ d[6] ^ c[30] ^ d[1] ^ d[10] ^ d[14] ^ d[5] ^ c[26] ^ c[18] ^ c[21] ^ d[18] ^ c[13] ^ c[25] ^ d[13] ;
o[22] = d[23] ^ c[17] ^ c[27] ^ c[20] ^ c[19] ^ c[22] ^ c[24] ^ d[12] ^ d[5] ^ c[26] ^ d[14] ^ c[8] ^ d[7] ^ d[0] ^ c[31] ^ d[9] ^ d[11] ^ d[4] ;
o[23] = d[23] ^ c[17] ^ c[27] ^ d[6] ^ c[9] ^ d[17] ^ d[8] ^ d[10] ^ c[14] ^ c[24] ^ d[3] ^ d[22] ^ d[14] ^ c[8] ^ d[7] ^ c[28] ^ c[21] ^ c[23] ^ d[4] ^ c[25] ;
o[24] = c[0] ^ d[6] ^ c[9] ^ c[10] ^ c[29] ^ c[22] ^ c[24] ^ d[3] ^ d[22] ^ d[5] ^ c[26] ^ c[18] ^ d[16] ^ d[7] ^ c[28] ^ d[9] ^ d[2] ^ c[15] ^ d[21] ^ c[25] ^ d[13] ;
o[25] = d[15] ^ d[6] ^ c[10] ^ c[27] ^ c[19] ^ c[29] ^ c[30] ^ d[8] ^ d[1] ^ d[20] ^ d[12] ^ c[16] ^ d[5] ^ c[26] ^ c[1] ^ c[11] ^ d[2] ^ c[23] ^ d[21] ^ c[25] ^ d[4] ;
o[26] = d[23] ^ c[27] ^ c[2] ^ d[17] ^ c[30] ^ c[12] ^ d[1] ^ c[14] ^ d[20] ^ d[19] ^ d[3] ^ d[5] ^ c[26] ^ c[8] ^ c[18] ^ c[28] ^ c[11] ^ d[0] ^ c[31] ^ d[4] ^ d[13] ;
o[27] = c[27] ^ c[9] ^ c[19] ^ c[29] ^ c[12] ^ d[19] ^ d[3] ^ d[12] ^ d[22] ^ d[16] ^ c[28] ^ d[0] ^ c[3] ^ c[31] ^ d[18] ^ c[13] ^ d[2] ^ c[15] ^ d[4] ;
o[28] = d[15] ^ c[10] ^ c[20] ^ c[29] ^ c[30] ^ d[17] ^ d[1] ^ c[4] ^ c[14] ^ d[3] ^ c[16] ^ c[28] ^ d[18] ^ c[13] ^ d[2] ^ d[11] ^ d[21] ;
o[29] = c[17] ^ c[29] ^ c[30] ^ d[17] ^ d[1] ^ d[10] ^ d[20] ^ c[14] ^ d[14] ^ c[11] ^ d[16] ^ d[0] ^ c[21] ^ c[31] ^ d[2] ^ c[5] ^ c[15] ;
o[30] = d[15] ^ c[30] ^ c[12] ^ d[1] ^ c[22] ^ d[19] ^ c[6] ^ c[16] ^ c[18] ^ d[16] ^ d[0] ^ c[31] ^ d[9] ^ c[15] ^ d[13] ;
o[31] = c[17] ^ d[15] ^ c[19] ^ d[8] ^ d[12] ^ c[16] ^ d[14] ^ d[0] ^ d[18] ^ c[31] ^ c[13] ^ c[23] ^ c[7] ;
        crc3B = o;
    end
    endfunction // crc3B

    ////////////////////////////////////////////////
    // crc2B
    ////////////////////////////////////////////////
    function [31:0] crc2B (
        input        [31:0]      c,
        input        [15:0]      d
        );
    reg          [31:0]      o;
    begin
o[0] = d[9] ^ c[22] ^ d[5] ^ c[26] ^ d[15] ^ d[6] ^ d[3] ^ c[28] ^ c[25] ^ c[16] ;
o[1] = c[17] ^ d[15] ^ d[6] ^ c[27] ^ c[29] ^ d[8] ^ c[22] ^ d[3] ^ c[16] ^ d[14] ^ c[28] ^ d[9] ^ c[23] ^ d[2] ^ d[4] ^ c[25] ;
o[2] = c[17] ^ d[15] ^ d[6] ^ d[8] ^ c[29] ^ c[30] ^ c[22] ^ d[1] ^ c[24] ^ c[16] ^ d[14] ^ c[18] ^ d[7] ^ d[9] ^ d[2] ^ c[23] ^ c[25] ^ d[13] ;
o[3] = c[17] ^ d[6] ^ c[19] ^ d[8] ^ c[30] ^ d[1] ^ c[24] ^ d[12] ^ d[14] ^ d[5] ^ c[26] ^ c[18] ^ d[7] ^ d[0] ^ c[31] ^ c[23] ^ d[13] ^ c[25] ;
o[4] = d[15] ^ c[27] ^ c[20] ^ c[19] ^ c[22] ^ d[3] ^ c[24] ^ d[12] ^ c[16] ^ c[18] ^ c[28] ^ d[7] ^ d[0] ^ d[9] ^ c[31] ^ d[11] ^ d[13] ^ d[4] ;
o[5] = c[17] ^ d[15] ^ c[19] ^ c[20] ^ d[8] ^ c[29] ^ c[22] ^ d[10] ^ d[12] ^ c[16] ^ d[5] ^ c[26] ^ d[14] ^ c[21] ^ d[9] ^ d[2] ^ c[23] ^ d[11] ;
o[6] = c[17] ^ c[27] ^ c[20] ^ d[8] ^ c[30] ^ d[1] ^ c[22] ^ d[10] ^ c[24] ^ d[14] ^ c[18] ^ d[7] ^ c[21] ^ d[9] ^ c[23] ^ d[11] ^ d[4] ^ d[13] ;
o[7] = d[15] ^ c[19] ^ d[8] ^ d[10] ^ c[24] ^ d[12] ^ c[16] ^ d[5] ^ c[26] ^ c[18] ^ d[7] ^ d[0] ^ c[21] ^ c[31] ^ c[23] ^ d[13] ;
o[8] = c[17] ^ d[15] ^ c[27] ^ c[19] ^ c[20] ^ d[3] ^ d[12] ^ c[24] ^ c[16] ^ d[5] ^ c[26] ^ d[14] ^ c[28] ^ d[7] ^ d[11] ^ d[4] ;
o[9] = c[17] ^ c[27] ^ d[6] ^ c[20] ^ c[29] ^ d[10] ^ d[3] ^ d[14] ^ c[18] ^ c[28] ^ c[21] ^ d[2] ^ d[11] ^ d[4] ^ d[13] ^ c[25] ;
o[10] = d[15] ^ d[6] ^ c[19] ^ c[30] ^ c[29] ^ d[1] ^ d[10] ^ d[12] ^ c[16] ^ c[18] ^ c[21] ^ d[2] ^ c[25] ^ d[13] ;
o[11] = c[17] ^ d[15] ^ d[6] ^ c[19] ^ c[20] ^ c[30] ^ d[1] ^ d[3] ^ d[12] ^ c[16] ^ d[14] ^ c[28] ^ d[0] ^ c[31] ^ d[11] ^ c[25] ;
o[12] = c[17] ^ d[15] ^ d[6] ^ c[20] ^ c[29] ^ c[22] ^ d[10] ^ d[3] ^ c[16] ^ d[14] ^ c[18] ^ c[28] ^ d[0] ^ c[21] ^ d[9] ^ c[31] ^ d[2] ^ d[11] ^ c[25] ^ d[13] ;
o[13] = c[17] ^ c[19] ^ d[8] ^ c[29] ^ c[30] ^ d[1] ^ d[10] ^ c[22] ^ d[12] ^ d[14] ^ d[5] ^ c[26] ^ c[18] ^ c[21] ^ d[9] ^ d[2] ^ c[23] ^ d[13] ;
o[14] = c[27] ^ c[19] ^ c[20] ^ c[30] ^ d[8] ^ d[1] ^ c[22] ^ c[24] ^ d[12] ^ c[18] ^ d[7] ^ d[0] ^ c[31] ^ d[9] ^ d[11] ^ c[23] ^ d[13] ^ d[4] ;
o[15] = d[6] ^ c[20] ^ c[19] ^ d[8] ^ d[10] ^ d[12] ^ c[24] ^ d[3] ^ d[7] ^ c[28] ^ d[0] ^ c[21] ^ c[31] ^ c[23] ^ d[11] ^ c[25] ;
o[16] = c[0] ^ d[15] ^ c[20] ^ c[29] ^ d[10] ^ d[3] ^ c[24] ^ c[16] ^ c[28] ^ d[7] ^ c[21] ^ d[11] ^ d[2] ;
o[17] = c[17] ^ d[6] ^ c[29] ^ c[30] ^ d[10] ^ d[1] ^ c[22] ^ d[14] ^ c[1] ^ c[21] ^ d[9] ^ d[2] ^ c[25] ;
o[18] = c[2] ^ c[30] ^ d[8] ^ d[1] ^ c[22] ^ c[26] ^ d[5] ^ c[18] ^ d[0] ^ d[9] ^ c[31] ^ c[23] ^ d[13] ;
o[19] = c[27] ^ c[19] ^ d[8] ^ d[12] ^ c[24] ^ d[7] ^ d[0] ^ c[3] ^ c[31] ^ c[23] ^ d[4] ;
o[20] = d[6] ^ c[20] ^ c[4] ^ d[3] ^ c[24] ^ d[7] ^ c[28] ^ d[11] ^ c[25] ;
o[21] = d[6] ^ c[29] ^ d[10] ^ c[26] ^ d[5] ^ c[21] ^ c[5] ^ d[2] ^ c[25] ;
o[22] = d[15] ^ d[6] ^ c[27] ^ c[30] ^ d[1] ^ d[3] ^ c[6] ^ c[16] ^ c[28] ^ c[25] ^ d[4] ;
o[23] = c[17] ^ d[15] ^ d[6] ^ c[29] ^ c[22] ^ c[16] ^ d[14] ^ d[0] ^ d[9] ^ c[31] ^ d[2] ^ c[25] ^ c[7] ;
o[24] = d[14] ^ d[5] ^ c[26] ^ c[17] ^ d[1] ^ c[8] ^ c[23] ^ c[18] ^ d[8] ^ d[13] ^ c[30] ;
o[25] = c[31] ^ c[27] ^ c[18] ^ c[9] ^ d[7] ^ c[24] ^ d[12] ^ c[19] ^ d[13] ^ d[4] ^ d[0] ;
o[26] = d[15] ^ c[10] ^ c[20] ^ c[19] ^ c[22] ^ d[12] ^ c[16] ^ d[5] ^ c[26] ^ d[9] ^ d[11] ;
o[27] = c[17] ^ c[27] ^ c[20] ^ d[8] ^ d[10] ^ d[14] ^ c[11] ^ c[21] ^ c[23] ^ d[11] ^ d[4] ;
o[28] = c[12] ^ c[22] ^ d[10] ^ c[24] ^ d[3] ^ c[18] ^ d[7] ^ c[28] ^ c[21] ^ d[9] ^ d[13] ;
o[29] = d[6] ^ c[19] ^ d[8] ^ c[29] ^ c[22] ^ d[12] ^ c[13] ^ d[9] ^ d[2] ^ c[23] ^ c[25] ;
o[30] = d[5] ^ c[26] ^ d[1] ^ d[11] ^ c[23] ^ c[14] ^ c[20] ^ d[7] ^ c[24] ^ c[30] ^ d[8] ;
o[31] = d[10] ^ c[31] ^ c[27] ^ d[6] ^ d[7] ^ c[24] ^ c[15] ^ d[4] ^ d[0] ^ c[21] ^ c[25] ;
        crc2B = o;
    end
    endfunction // crc2B

    ////////////////////////////////////////////////
    // crc1B
    ////////////////////////////////////////////////
    function [31:0] crc1B (
        input        [31:0]      c,
        input        [7:0]       d
        );
    reg          [31:0]      o;
    begin
o[0] = d[1] ^ d[7] ^ c[24] ^ c[30] ;
o[1] = d[1] ^ c[31] ^ d[6] ^ d[7] ^ c[24] ^ c[30] ^ d[0] ^ c[25] ;
o[2] = d[1] ^ c[31] ^ d[5] ^ c[26] ^ d[6] ^ d[7] ^ c[24] ^ c[30] ^ d[0] ^ c[25] ;
o[3] = c[31] ^ d[5] ^ c[26] ^ d[6] ^ c[27] ^ d[0] ^ c[25] ^ d[4] ;
o[4] = d[1] ^ d[5] ^ c[26] ^ c[27] ^ d[7] ^ c[24] ^ d[3] ^ c[28] ^ c[30] ^ d[4] ;
o[5] = c[27] ^ d[6] ^ c[30] ^ c[29] ^ d[1] ^ d[3] ^ c[24] ^ d[7] ^ c[28] ^ d[0] ^ c[31] ^ d[2] ^ d[4] ^ c[25] ;
o[6] = d[6] ^ c[30] ^ c[29] ^ d[1] ^ d[3] ^ c[26] ^ d[5] ^ c[28] ^ d[0] ^ c[31] ^ d[2] ^ c[25] ;
o[7] = d[5] ^ c[26] ^ c[31] ^ c[27] ^ d[2] ^ d[7] ^ c[24] ^ d[4] ^ c[29] ^ d[0] ;
o[8] = c[0] ^ d[6] ^ c[27] ^ d[7] ^ c[24] ^ d[3] ^ c[28] ^ c[25] ^ d[4] ;
o[9] = d[5] ^ c[26] ^ d[6] ^ d[2] ^ c[1] ^ d[3] ^ c[28] ^ c[25] ^ c[29] ;
o[10] = d[5] ^ c[26] ^ c[27] ^ d[2] ^ d[7] ^ c[24] ^ c[2] ^ d[4] ^ c[29] ;
o[11] = d[6] ^ c[27] ^ d[7] ^ c[24] ^ d[3] ^ c[28] ^ c[25] ^ d[4] ^ c[3] ;
o[12] = d[6] ^ c[29] ^ c[30] ^ d[1] ^ c[4] ^ d[3] ^ c[24] ^ c[26] ^ d[5] ^ d[7] ^ c[28] ^ d[2] ^ c[25] ;
o[13] = d[6] ^ c[27] ^ c[30] ^ c[29] ^ d[1] ^ c[26] ^ d[5] ^ d[0] ^ c[31] ^ c[5] ^ d[2] ^ d[4] ^ c[25] ;
o[14] = d[5] ^ c[26] ^ d[1] ^ c[31] ^ c[27] ^ d[3] ^ c[28] ^ c[6] ^ d[4] ^ c[30] ^ d[0] ;
o[15] = c[31] ^ c[27] ^ d[2] ^ d[3] ^ c[28] ^ d[4] ^ c[29] ^ d[0] ^ c[7] ;
o[16] = c[8] ^ d[2] ^ d[7] ^ c[24] ^ d[3] ^ c[28] ^ c[29] ;
o[17] = d[1] ^ d[6] ^ d[2] ^ c[9] ^ c[25] ^ c[29] ^ c[30] ;
o[18] = d[5] ^ c[26] ^ d[1] ^ c[31] ^ c[10] ^ c[30] ^ d[0] ;
o[19] = c[31] ^ c[27] ^ c[11] ^ d[4] ^ d[0] ;
o[20] = d[3] ^ c[28] ^ c[12] ;
o[21] = c[13] ^ d[2] ^ c[29] ;
o[22] = c[14] ^ d[7] ^ c[24] ;
o[23] = d[1] ^ d[6] ^ d[7] ^ c[24] ^ c[15] ^ c[30] ^ c[25] ;
o[24] = c[31] ^ d[5] ^ c[26] ^ d[6] ^ d[0] ^ c[25] ^ c[16] ;
o[25] = d[5] ^ c[26] ^ c[17] ^ c[27] ^ d[4] ;
o[26] = d[1] ^ c[27] ^ c[18] ^ d[7] ^ c[24] ^ d[3] ^ c[28] ^ c[30] ^ d[4] ;
o[27] = c[31] ^ d[6] ^ d[2] ^ d[3] ^ c[28] ^ c[19] ^ d[0] ^ c[25] ^ c[29] ;
o[28] = d[5] ^ c[26] ^ d[1] ^ d[2] ^ c[20] ^ c[29] ^ c[30] ;
o[29] = d[1] ^ c[31] ^ c[27] ^ d[4] ^ c[30] ^ d[0] ^ c[21] ;
o[30] = c[31] ^ c[22] ^ d[3] ^ c[28] ^ d[0] ;
o[31] = d[2] ^ c[23] ^ c[29] ;
        crc1B = o;
    end
    endfunction // crc1B

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////